
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"e8",x"d2",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"e8",x"d2",x"c2"),
    14 => (x"48",x"f4",x"c0",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"c8",x"ff"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d6",x"02",x"99"),
    50 => (x"c3",x"48",x"d4",x"ff"),
    51 => (x"52",x"68",x"78",x"ff"),
    52 => (x"48",x"49",x"66",x"c4"),
    53 => (x"a6",x"c8",x"88",x"c1"),
    54 => (x"05",x"99",x"71",x"58"),
    55 => (x"4f",x"26",x"87",x"ea"),
    56 => (x"ff",x"1e",x"73",x"1e"),
    57 => (x"ff",x"c3",x"4b",x"d4"),
    58 => (x"c3",x"4a",x"6b",x"7b"),
    59 => (x"49",x"6b",x"7b",x"ff"),
    60 => (x"b1",x"72",x"32",x"c8"),
    61 => (x"6b",x"7b",x"ff",x"c3"),
    62 => (x"71",x"31",x"c8",x"4a"),
    63 => (x"7b",x"ff",x"c3",x"b2"),
    64 => (x"32",x"c8",x"49",x"6b"),
    65 => (x"48",x"71",x"b1",x"72"),
    66 => (x"4d",x"26",x"87",x"c4"),
    67 => (x"4b",x"26",x"4c",x"26"),
    68 => (x"5e",x"0e",x"4f",x"26"),
    69 => (x"0e",x"5d",x"5c",x"5b"),
    70 => (x"d4",x"ff",x"4a",x"71"),
    71 => (x"c3",x"49",x"72",x"4c"),
    72 => (x"7c",x"71",x"99",x"ff"),
    73 => (x"bf",x"f4",x"c0",x"c2"),
    74 => (x"d0",x"87",x"c8",x"05"),
    75 => (x"30",x"c9",x"48",x"66"),
    76 => (x"d0",x"58",x"a6",x"d4"),
    77 => (x"29",x"d8",x"49",x"66"),
    78 => (x"71",x"99",x"ff",x"c3"),
    79 => (x"49",x"66",x"d0",x"7c"),
    80 => (x"ff",x"c3",x"29",x"d0"),
    81 => (x"d0",x"7c",x"71",x"99"),
    82 => (x"29",x"c8",x"49",x"66"),
    83 => (x"71",x"99",x"ff",x"c3"),
    84 => (x"49",x"66",x"d0",x"7c"),
    85 => (x"71",x"99",x"ff",x"c3"),
    86 => (x"d0",x"49",x"72",x"7c"),
    87 => (x"99",x"ff",x"c3",x"29"),
    88 => (x"4b",x"6c",x"7c",x"71"),
    89 => (x"4d",x"ff",x"f0",x"c9"),
    90 => (x"05",x"ab",x"ff",x"c3"),
    91 => (x"ff",x"c3",x"87",x"d0"),
    92 => (x"c1",x"4b",x"6c",x"7c"),
    93 => (x"87",x"c6",x"02",x"8d"),
    94 => (x"02",x"ab",x"ff",x"c3"),
    95 => (x"48",x"73",x"87",x"f0"),
    96 => (x"0e",x"87",x"c7",x"fe"),
    97 => (x"5d",x"5c",x"5b",x"5e"),
    98 => (x"c0",x"4b",x"71",x"0e"),
    99 => (x"cd",x"ee",x"c5",x"4c"),
   100 => (x"d4",x"ff",x"4a",x"df"),
   101 => (x"78",x"ff",x"c3",x"48"),
   102 => (x"fe",x"c3",x"49",x"68"),
   103 => (x"fd",x"c0",x"05",x"a9"),
   104 => (x"73",x"4d",x"70",x"87"),
   105 => (x"87",x"cc",x"02",x"9b"),
   106 => (x"73",x"1e",x"66",x"d0"),
   107 => (x"87",x"c7",x"fc",x"49"),
   108 => (x"87",x"d6",x"86",x"c4"),
   109 => (x"c4",x"48",x"d0",x"ff"),
   110 => (x"ff",x"c3",x"78",x"d1"),
   111 => (x"48",x"66",x"d0",x"7d"),
   112 => (x"a6",x"d4",x"88",x"c1"),
   113 => (x"05",x"98",x"70",x"58"),
   114 => (x"d4",x"ff",x"87",x"f0"),
   115 => (x"78",x"ff",x"c3",x"48"),
   116 => (x"05",x"9b",x"73",x"78"),
   117 => (x"d0",x"ff",x"87",x"c5"),
   118 => (x"c1",x"78",x"d0",x"48"),
   119 => (x"8a",x"c1",x"4c",x"4a"),
   120 => (x"87",x"ee",x"fe",x"05"),
   121 => (x"e1",x"fc",x"48",x"74"),
   122 => (x"1e",x"73",x"1e",x"87"),
   123 => (x"4b",x"c0",x"4a",x"71"),
   124 => (x"c3",x"48",x"d4",x"ff"),
   125 => (x"d0",x"ff",x"78",x"ff"),
   126 => (x"78",x"c3",x"c4",x"48"),
   127 => (x"c3",x"48",x"d4",x"ff"),
   128 => (x"1e",x"72",x"78",x"ff"),
   129 => (x"c1",x"f0",x"ff",x"c0"),
   130 => (x"c5",x"fc",x"49",x"d1"),
   131 => (x"70",x"86",x"c4",x"87"),
   132 => (x"87",x"d2",x"05",x"98"),
   133 => (x"cc",x"1e",x"c0",x"c8"),
   134 => (x"e6",x"fd",x"49",x"66"),
   135 => (x"70",x"86",x"c4",x"87"),
   136 => (x"48",x"d0",x"ff",x"4b"),
   137 => (x"48",x"73",x"78",x"c2"),
   138 => (x"0e",x"87",x"e3",x"fb"),
   139 => (x"5d",x"5c",x"5b",x"5e"),
   140 => (x"c2",x"86",x"f8",x"0e"),
   141 => (x"c0",x"48",x"cc",x"c9"),
   142 => (x"c4",x"c1",x"c2",x"78"),
   143 => (x"fe",x"49",x"c0",x"1e"),
   144 => (x"86",x"c4",x"87",x"e7"),
   145 => (x"c5",x"05",x"98",x"70"),
   146 => (x"c9",x"48",x"c0",x"87"),
   147 => (x"4d",x"c0",x"87",x"cc"),
   148 => (x"e4",x"c0",x"7e",x"c1"),
   149 => (x"c2",x"49",x"bf",x"cf"),
   150 => (x"71",x"4a",x"fa",x"c1"),
   151 => (x"c8",x"f8",x"4b",x"c8"),
   152 => (x"05",x"98",x"70",x"87"),
   153 => (x"7e",x"c0",x"87",x"c2"),
   154 => (x"bf",x"cb",x"e4",x"c0"),
   155 => (x"d6",x"c2",x"c2",x"49"),
   156 => (x"4b",x"c8",x"71",x"4a"),
   157 => (x"70",x"87",x"f2",x"f7"),
   158 => (x"87",x"c2",x"05",x"98"),
   159 => (x"02",x"6e",x"7e",x"c0"),
   160 => (x"c2",x"87",x"fd",x"c0"),
   161 => (x"4d",x"bf",x"ca",x"c8"),
   162 => (x"9f",x"c2",x"c9",x"c2"),
   163 => (x"c5",x"48",x"7e",x"bf"),
   164 => (x"05",x"a8",x"ea",x"d6"),
   165 => (x"c8",x"c2",x"87",x"c7"),
   166 => (x"ce",x"4d",x"bf",x"ca"),
   167 => (x"ca",x"48",x"6e",x"87"),
   168 => (x"02",x"a8",x"d5",x"e9"),
   169 => (x"48",x"c0",x"87",x"c5"),
   170 => (x"c2",x"87",x"ef",x"c7"),
   171 => (x"75",x"1e",x"c4",x"c1"),
   172 => (x"87",x"f5",x"fc",x"49"),
   173 => (x"98",x"70",x"86",x"c4"),
   174 => (x"c0",x"87",x"c5",x"05"),
   175 => (x"87",x"da",x"c7",x"48"),
   176 => (x"bf",x"cb",x"e4",x"c0"),
   177 => (x"d6",x"c2",x"c2",x"49"),
   178 => (x"4b",x"c8",x"71",x"4a"),
   179 => (x"70",x"87",x"da",x"f6"),
   180 => (x"87",x"c8",x"05",x"98"),
   181 => (x"48",x"cc",x"c9",x"c2"),
   182 => (x"87",x"d9",x"78",x"c1"),
   183 => (x"bf",x"cf",x"e4",x"c0"),
   184 => (x"fa",x"c1",x"c2",x"49"),
   185 => (x"4b",x"c8",x"71",x"4a"),
   186 => (x"70",x"87",x"fe",x"f5"),
   187 => (x"87",x"c5",x"02",x"98"),
   188 => (x"e5",x"c6",x"48",x"c0"),
   189 => (x"c2",x"c9",x"c2",x"87"),
   190 => (x"c1",x"49",x"bf",x"97"),
   191 => (x"cd",x"05",x"a9",x"d5"),
   192 => (x"c3",x"c9",x"c2",x"87"),
   193 => (x"c2",x"49",x"bf",x"97"),
   194 => (x"c0",x"02",x"a9",x"ea"),
   195 => (x"48",x"c0",x"87",x"c5"),
   196 => (x"c2",x"87",x"c7",x"c6"),
   197 => (x"bf",x"97",x"c4",x"c1"),
   198 => (x"e9",x"c3",x"48",x"7e"),
   199 => (x"ce",x"c0",x"02",x"a8"),
   200 => (x"c3",x"48",x"6e",x"87"),
   201 => (x"c0",x"02",x"a8",x"eb"),
   202 => (x"48",x"c0",x"87",x"c5"),
   203 => (x"c2",x"87",x"eb",x"c5"),
   204 => (x"bf",x"97",x"cf",x"c1"),
   205 => (x"c0",x"05",x"99",x"49"),
   206 => (x"c1",x"c2",x"87",x"cc"),
   207 => (x"49",x"bf",x"97",x"d0"),
   208 => (x"c0",x"02",x"a9",x"c2"),
   209 => (x"48",x"c0",x"87",x"c5"),
   210 => (x"c2",x"87",x"cf",x"c5"),
   211 => (x"bf",x"97",x"d1",x"c1"),
   212 => (x"c8",x"c9",x"c2",x"48"),
   213 => (x"48",x"4c",x"70",x"58"),
   214 => (x"c9",x"c2",x"88",x"c1"),
   215 => (x"c1",x"c2",x"58",x"cc"),
   216 => (x"49",x"bf",x"97",x"d2"),
   217 => (x"c1",x"c2",x"81",x"75"),
   218 => (x"4a",x"bf",x"97",x"d3"),
   219 => (x"a1",x"72",x"32",x"c8"),
   220 => (x"d9",x"cd",x"c2",x"7e"),
   221 => (x"c2",x"78",x"6e",x"48"),
   222 => (x"bf",x"97",x"d4",x"c1"),
   223 => (x"58",x"a6",x"c8",x"48"),
   224 => (x"bf",x"cc",x"c9",x"c2"),
   225 => (x"87",x"d4",x"c2",x"02"),
   226 => (x"bf",x"cb",x"e4",x"c0"),
   227 => (x"d6",x"c2",x"c2",x"49"),
   228 => (x"4b",x"c8",x"71",x"4a"),
   229 => (x"70",x"87",x"d2",x"f3"),
   230 => (x"c5",x"c0",x"02",x"98"),
   231 => (x"c3",x"48",x"c0",x"87"),
   232 => (x"c9",x"c2",x"87",x"f8"),
   233 => (x"c2",x"4c",x"bf",x"c4"),
   234 => (x"c2",x"5c",x"ed",x"cd"),
   235 => (x"bf",x"97",x"e9",x"c1"),
   236 => (x"c2",x"31",x"c8",x"49"),
   237 => (x"bf",x"97",x"e8",x"c1"),
   238 => (x"c2",x"49",x"a1",x"4a"),
   239 => (x"bf",x"97",x"ea",x"c1"),
   240 => (x"72",x"32",x"d0",x"4a"),
   241 => (x"c1",x"c2",x"49",x"a1"),
   242 => (x"4a",x"bf",x"97",x"eb"),
   243 => (x"a1",x"72",x"32",x"d8"),
   244 => (x"91",x"66",x"c4",x"49"),
   245 => (x"bf",x"d9",x"cd",x"c2"),
   246 => (x"e1",x"cd",x"c2",x"81"),
   247 => (x"f1",x"c1",x"c2",x"59"),
   248 => (x"c8",x"4a",x"bf",x"97"),
   249 => (x"f0",x"c1",x"c2",x"32"),
   250 => (x"a2",x"4b",x"bf",x"97"),
   251 => (x"f2",x"c1",x"c2",x"4a"),
   252 => (x"d0",x"4b",x"bf",x"97"),
   253 => (x"4a",x"a2",x"73",x"33"),
   254 => (x"97",x"f3",x"c1",x"c2"),
   255 => (x"9b",x"cf",x"4b",x"bf"),
   256 => (x"a2",x"73",x"33",x"d8"),
   257 => (x"e5",x"cd",x"c2",x"4a"),
   258 => (x"e1",x"cd",x"c2",x"5a"),
   259 => (x"8a",x"c2",x"4a",x"bf"),
   260 => (x"cd",x"c2",x"92",x"74"),
   261 => (x"a1",x"72",x"48",x"e5"),
   262 => (x"87",x"ca",x"c1",x"78"),
   263 => (x"97",x"d6",x"c1",x"c2"),
   264 => (x"31",x"c8",x"49",x"bf"),
   265 => (x"97",x"d5",x"c1",x"c2"),
   266 => (x"49",x"a1",x"4a",x"bf"),
   267 => (x"59",x"d4",x"c9",x"c2"),
   268 => (x"bf",x"d0",x"c9",x"c2"),
   269 => (x"c7",x"31",x"c5",x"49"),
   270 => (x"29",x"c9",x"81",x"ff"),
   271 => (x"59",x"ed",x"cd",x"c2"),
   272 => (x"97",x"db",x"c1",x"c2"),
   273 => (x"32",x"c8",x"4a",x"bf"),
   274 => (x"97",x"da",x"c1",x"c2"),
   275 => (x"4a",x"a2",x"4b",x"bf"),
   276 => (x"6e",x"92",x"66",x"c4"),
   277 => (x"e9",x"cd",x"c2",x"82"),
   278 => (x"e1",x"cd",x"c2",x"5a"),
   279 => (x"c2",x"78",x"c0",x"48"),
   280 => (x"72",x"48",x"dd",x"cd"),
   281 => (x"cd",x"c2",x"78",x"a1"),
   282 => (x"cd",x"c2",x"48",x"ed"),
   283 => (x"c2",x"78",x"bf",x"e1"),
   284 => (x"c2",x"48",x"f1",x"cd"),
   285 => (x"78",x"bf",x"e5",x"cd"),
   286 => (x"bf",x"cc",x"c9",x"c2"),
   287 => (x"87",x"c9",x"c0",x"02"),
   288 => (x"30",x"c4",x"48",x"74"),
   289 => (x"c9",x"c0",x"7e",x"70"),
   290 => (x"e9",x"cd",x"c2",x"87"),
   291 => (x"30",x"c4",x"48",x"bf"),
   292 => (x"c9",x"c2",x"7e",x"70"),
   293 => (x"78",x"6e",x"48",x"d0"),
   294 => (x"8e",x"f8",x"48",x"c1"),
   295 => (x"4c",x"26",x"4d",x"26"),
   296 => (x"4f",x"26",x"4b",x"26"),
   297 => (x"5c",x"5b",x"5e",x"0e"),
   298 => (x"4a",x"71",x"0e",x"5d"),
   299 => (x"bf",x"cc",x"c9",x"c2"),
   300 => (x"72",x"87",x"cb",x"02"),
   301 => (x"72",x"2b",x"c7",x"4b"),
   302 => (x"9c",x"ff",x"c1",x"4c"),
   303 => (x"4b",x"72",x"87",x"c9"),
   304 => (x"4c",x"72",x"2b",x"c8"),
   305 => (x"c2",x"9c",x"ff",x"c3"),
   306 => (x"83",x"bf",x"d9",x"cd"),
   307 => (x"bf",x"c7",x"e4",x"c0"),
   308 => (x"87",x"d9",x"02",x"ab"),
   309 => (x"5b",x"cb",x"e4",x"c0"),
   310 => (x"1e",x"c4",x"c1",x"c2"),
   311 => (x"c8",x"f4",x"49",x"73"),
   312 => (x"70",x"86",x"c4",x"87"),
   313 => (x"87",x"c5",x"05",x"98"),
   314 => (x"e6",x"c0",x"48",x"c0"),
   315 => (x"cc",x"c9",x"c2",x"87"),
   316 => (x"87",x"d2",x"02",x"bf"),
   317 => (x"91",x"c4",x"49",x"74"),
   318 => (x"81",x"c4",x"c1",x"c2"),
   319 => (x"ff",x"cf",x"4d",x"69"),
   320 => (x"9d",x"ff",x"ff",x"ff"),
   321 => (x"49",x"74",x"87",x"cb"),
   322 => (x"c1",x"c2",x"91",x"c2"),
   323 => (x"69",x"9f",x"81",x"c4"),
   324 => (x"fe",x"48",x"75",x"4d"),
   325 => (x"5e",x"0e",x"87",x"c6"),
   326 => (x"0e",x"5d",x"5c",x"5b"),
   327 => (x"4c",x"71",x"86",x"f8"),
   328 => (x"87",x"c5",x"05",x"9c"),
   329 => (x"c1",x"c3",x"48",x"c0"),
   330 => (x"7e",x"a4",x"c8",x"87"),
   331 => (x"d8",x"78",x"c0",x"48"),
   332 => (x"87",x"c7",x"02",x"66"),
   333 => (x"bf",x"97",x"66",x"d8"),
   334 => (x"c0",x"87",x"c5",x"05"),
   335 => (x"87",x"ea",x"c2",x"48"),
   336 => (x"49",x"c1",x"1e",x"c0"),
   337 => (x"87",x"e6",x"c7",x"49"),
   338 => (x"4d",x"70",x"86",x"c4"),
   339 => (x"c2",x"c1",x"02",x"9d"),
   340 => (x"d4",x"c9",x"c2",x"87"),
   341 => (x"49",x"66",x"d8",x"4a"),
   342 => (x"70",x"87",x"f3",x"eb"),
   343 => (x"f2",x"c0",x"02",x"98"),
   344 => (x"d8",x"4a",x"75",x"87"),
   345 => (x"4b",x"cb",x"49",x"66"),
   346 => (x"70",x"87",x"d8",x"ec"),
   347 => (x"e2",x"c0",x"02",x"98"),
   348 => (x"75",x"1e",x"c0",x"87"),
   349 => (x"87",x"c7",x"02",x"9d"),
   350 => (x"c0",x"48",x"a6",x"c8"),
   351 => (x"c8",x"87",x"c5",x"78"),
   352 => (x"78",x"c1",x"48",x"a6"),
   353 => (x"c6",x"49",x"66",x"c8"),
   354 => (x"86",x"c4",x"87",x"e4"),
   355 => (x"05",x"9d",x"4d",x"70"),
   356 => (x"75",x"87",x"fe",x"fe"),
   357 => (x"cf",x"c1",x"02",x"9d"),
   358 => (x"49",x"a5",x"dc",x"87"),
   359 => (x"78",x"69",x"48",x"6e"),
   360 => (x"c4",x"49",x"a5",x"da"),
   361 => (x"a4",x"c4",x"48",x"a6"),
   362 => (x"48",x"69",x"9f",x"78"),
   363 => (x"78",x"08",x"66",x"c4"),
   364 => (x"bf",x"cc",x"c9",x"c2"),
   365 => (x"d4",x"87",x"d2",x"02"),
   366 => (x"69",x"9f",x"49",x"a5"),
   367 => (x"ff",x"ff",x"c0",x"49"),
   368 => (x"d0",x"48",x"71",x"99"),
   369 => (x"c2",x"7e",x"70",x"30"),
   370 => (x"6e",x"7e",x"c0",x"87"),
   371 => (x"66",x"c4",x"48",x"49"),
   372 => (x"66",x"c4",x"80",x"bf"),
   373 => (x"7c",x"c0",x"78",x"08"),
   374 => (x"c4",x"49",x"a4",x"cc"),
   375 => (x"d0",x"79",x"bf",x"66"),
   376 => (x"79",x"c0",x"49",x"a4"),
   377 => (x"87",x"c2",x"48",x"c1"),
   378 => (x"8e",x"f8",x"48",x"c0"),
   379 => (x"0e",x"87",x"ed",x"fa"),
   380 => (x"5d",x"5c",x"5b",x"5e"),
   381 => (x"9c",x"4c",x"71",x"0e"),
   382 => (x"87",x"ca",x"c1",x"02"),
   383 => (x"69",x"49",x"a4",x"c8"),
   384 => (x"87",x"c2",x"c1",x"02"),
   385 => (x"6c",x"4a",x"66",x"d0"),
   386 => (x"a6",x"d4",x"82",x"49"),
   387 => (x"4d",x"66",x"d0",x"5a"),
   388 => (x"c8",x"c9",x"c2",x"b9"),
   389 => (x"ba",x"ff",x"4a",x"bf"),
   390 => (x"99",x"71",x"99",x"72"),
   391 => (x"87",x"e4",x"c0",x"02"),
   392 => (x"6b",x"4b",x"a4",x"c4"),
   393 => (x"87",x"fc",x"f9",x"49"),
   394 => (x"c9",x"c2",x"7b",x"70"),
   395 => (x"6c",x"49",x"bf",x"c4"),
   396 => (x"75",x"7c",x"71",x"81"),
   397 => (x"c8",x"c9",x"c2",x"b9"),
   398 => (x"ba",x"ff",x"4a",x"bf"),
   399 => (x"99",x"71",x"99",x"72"),
   400 => (x"87",x"dc",x"ff",x"05"),
   401 => (x"d3",x"f9",x"7c",x"75"),
   402 => (x"1e",x"73",x"1e",x"87"),
   403 => (x"02",x"9b",x"4b",x"71"),
   404 => (x"a3",x"c8",x"87",x"c7"),
   405 => (x"c5",x"05",x"69",x"49"),
   406 => (x"c0",x"48",x"c0",x"87"),
   407 => (x"cd",x"c2",x"87",x"f7"),
   408 => (x"c4",x"4a",x"bf",x"dd"),
   409 => (x"49",x"69",x"49",x"a3"),
   410 => (x"c9",x"c2",x"89",x"c2"),
   411 => (x"71",x"91",x"bf",x"c4"),
   412 => (x"c9",x"c2",x"4a",x"a2"),
   413 => (x"6b",x"49",x"bf",x"c8"),
   414 => (x"4a",x"a2",x"71",x"99"),
   415 => (x"5a",x"cb",x"e4",x"c0"),
   416 => (x"72",x"1e",x"66",x"c8"),
   417 => (x"87",x"e1",x"ed",x"49"),
   418 => (x"98",x"70",x"86",x"c4"),
   419 => (x"c0",x"87",x"c4",x"05"),
   420 => (x"c1",x"87",x"c2",x"48"),
   421 => (x"87",x"c8",x"f8",x"48"),
   422 => (x"71",x"1e",x"73",x"1e"),
   423 => (x"c0",x"02",x"9b",x"4b"),
   424 => (x"cd",x"c2",x"87",x"e4"),
   425 => (x"4a",x"73",x"5b",x"f1"),
   426 => (x"c9",x"c2",x"8a",x"c2"),
   427 => (x"92",x"49",x"bf",x"c4"),
   428 => (x"bf",x"dd",x"cd",x"c2"),
   429 => (x"c2",x"80",x"72",x"48"),
   430 => (x"71",x"58",x"f5",x"cd"),
   431 => (x"c2",x"30",x"c4",x"48"),
   432 => (x"c0",x"58",x"d4",x"c9"),
   433 => (x"cd",x"c2",x"87",x"ed"),
   434 => (x"cd",x"c2",x"48",x"ed"),
   435 => (x"c2",x"78",x"bf",x"e1"),
   436 => (x"c2",x"48",x"f1",x"cd"),
   437 => (x"78",x"bf",x"e5",x"cd"),
   438 => (x"bf",x"cc",x"c9",x"c2"),
   439 => (x"c2",x"87",x"c9",x"02"),
   440 => (x"49",x"bf",x"c4",x"c9"),
   441 => (x"87",x"c7",x"31",x"c4"),
   442 => (x"bf",x"e9",x"cd",x"c2"),
   443 => (x"c2",x"31",x"c4",x"49"),
   444 => (x"f6",x"59",x"d4",x"c9"),
   445 => (x"5e",x"0e",x"87",x"ea"),
   446 => (x"71",x"0e",x"5c",x"5b"),
   447 => (x"72",x"4b",x"c0",x"4a"),
   448 => (x"e1",x"c0",x"02",x"9a"),
   449 => (x"49",x"a2",x"da",x"87"),
   450 => (x"c2",x"4b",x"69",x"9f"),
   451 => (x"02",x"bf",x"cc",x"c9"),
   452 => (x"a2",x"d4",x"87",x"cf"),
   453 => (x"49",x"69",x"9f",x"49"),
   454 => (x"ff",x"ff",x"c0",x"4c"),
   455 => (x"c2",x"34",x"d0",x"9c"),
   456 => (x"74",x"4c",x"c0",x"87"),
   457 => (x"49",x"73",x"b3",x"49"),
   458 => (x"f5",x"87",x"ed",x"fd"),
   459 => (x"5e",x"0e",x"87",x"f0"),
   460 => (x"0e",x"5d",x"5c",x"5b"),
   461 => (x"4a",x"71",x"86",x"f4"),
   462 => (x"9a",x"72",x"7e",x"c0"),
   463 => (x"c2",x"87",x"d8",x"02"),
   464 => (x"c0",x"48",x"c0",x"c1"),
   465 => (x"f8",x"c0",x"c2",x"78"),
   466 => (x"f1",x"cd",x"c2",x"48"),
   467 => (x"c0",x"c2",x"78",x"bf"),
   468 => (x"cd",x"c2",x"48",x"fc"),
   469 => (x"c2",x"78",x"bf",x"ed"),
   470 => (x"c0",x"48",x"e1",x"c9"),
   471 => (x"d0",x"c9",x"c2",x"50"),
   472 => (x"c1",x"c2",x"49",x"bf"),
   473 => (x"71",x"4a",x"bf",x"c0"),
   474 => (x"c7",x"c4",x"03",x"aa"),
   475 => (x"cf",x"49",x"72",x"87"),
   476 => (x"e9",x"c0",x"05",x"99"),
   477 => (x"c7",x"e4",x"c0",x"87"),
   478 => (x"f8",x"c0",x"c2",x"48"),
   479 => (x"c1",x"c2",x"78",x"bf"),
   480 => (x"c0",x"c2",x"1e",x"c4"),
   481 => (x"c2",x"49",x"bf",x"f8"),
   482 => (x"c1",x"48",x"f8",x"c0"),
   483 => (x"e9",x"71",x"78",x"a1"),
   484 => (x"86",x"c4",x"87",x"d7"),
   485 => (x"48",x"c3",x"e4",x"c0"),
   486 => (x"78",x"c4",x"c1",x"c2"),
   487 => (x"e4",x"c0",x"87",x"cc"),
   488 => (x"c0",x"48",x"bf",x"c3"),
   489 => (x"e4",x"c0",x"80",x"e0"),
   490 => (x"c1",x"c2",x"58",x"c7"),
   491 => (x"c1",x"48",x"bf",x"c0"),
   492 => (x"c4",x"c1",x"c2",x"80"),
   493 => (x"09",x"03",x"27",x"58"),
   494 => (x"97",x"bf",x"00",x"00"),
   495 => (x"02",x"9d",x"4d",x"bf"),
   496 => (x"c3",x"87",x"e1",x"c2"),
   497 => (x"c2",x"02",x"ad",x"e5"),
   498 => (x"e4",x"c0",x"87",x"da"),
   499 => (x"cb",x"4b",x"bf",x"c3"),
   500 => (x"4c",x"11",x"49",x"a3"),
   501 => (x"c1",x"05",x"ac",x"cf"),
   502 => (x"49",x"75",x"87",x"d2"),
   503 => (x"89",x"c1",x"99",x"df"),
   504 => (x"c9",x"c2",x"91",x"cd"),
   505 => (x"a3",x"c1",x"81",x"d4"),
   506 => (x"c3",x"51",x"12",x"4a"),
   507 => (x"51",x"12",x"4a",x"a3"),
   508 => (x"12",x"4a",x"a3",x"c5"),
   509 => (x"4a",x"a3",x"c7",x"51"),
   510 => (x"a3",x"c9",x"51",x"12"),
   511 => (x"ce",x"51",x"12",x"4a"),
   512 => (x"51",x"12",x"4a",x"a3"),
   513 => (x"12",x"4a",x"a3",x"d0"),
   514 => (x"4a",x"a3",x"d2",x"51"),
   515 => (x"a3",x"d4",x"51",x"12"),
   516 => (x"d6",x"51",x"12",x"4a"),
   517 => (x"51",x"12",x"4a",x"a3"),
   518 => (x"12",x"4a",x"a3",x"d8"),
   519 => (x"4a",x"a3",x"dc",x"51"),
   520 => (x"a3",x"de",x"51",x"12"),
   521 => (x"c1",x"51",x"12",x"4a"),
   522 => (x"87",x"f8",x"c0",x"7e"),
   523 => (x"99",x"c8",x"49",x"74"),
   524 => (x"87",x"e9",x"c0",x"05"),
   525 => (x"99",x"d0",x"49",x"74"),
   526 => (x"dc",x"87",x"cf",x"05"),
   527 => (x"87",x"ca",x"02",x"66"),
   528 => (x"66",x"dc",x"49",x"73"),
   529 => (x"02",x"98",x"70",x"0f"),
   530 => (x"05",x"6e",x"87",x"d3"),
   531 => (x"c2",x"87",x"c6",x"c0"),
   532 => (x"c0",x"48",x"d4",x"c9"),
   533 => (x"c3",x"e4",x"c0",x"50"),
   534 => (x"e1",x"c2",x"48",x"bf"),
   535 => (x"e1",x"c9",x"c2",x"87"),
   536 => (x"7e",x"50",x"c0",x"48"),
   537 => (x"bf",x"d0",x"c9",x"c2"),
   538 => (x"c0",x"c1",x"c2",x"49"),
   539 => (x"aa",x"71",x"4a",x"bf"),
   540 => (x"87",x"f9",x"fb",x"04"),
   541 => (x"bf",x"f1",x"cd",x"c2"),
   542 => (x"87",x"c8",x"c0",x"05"),
   543 => (x"bf",x"cc",x"c9",x"c2"),
   544 => (x"87",x"f8",x"c1",x"02"),
   545 => (x"bf",x"fc",x"c0",x"c2"),
   546 => (x"87",x"d8",x"f0",x"49"),
   547 => (x"c1",x"c2",x"49",x"70"),
   548 => (x"a6",x"c4",x"59",x"c0"),
   549 => (x"fc",x"c0",x"c2",x"48"),
   550 => (x"c9",x"c2",x"78",x"bf"),
   551 => (x"c0",x"02",x"bf",x"cc"),
   552 => (x"66",x"c4",x"87",x"d8"),
   553 => (x"ff",x"ff",x"cf",x"49"),
   554 => (x"a9",x"99",x"f8",x"ff"),
   555 => (x"87",x"c5",x"c0",x"02"),
   556 => (x"e1",x"c0",x"4c",x"c0"),
   557 => (x"c0",x"4c",x"c1",x"87"),
   558 => (x"66",x"c4",x"87",x"dc"),
   559 => (x"f8",x"ff",x"cf",x"49"),
   560 => (x"c0",x"02",x"a9",x"99"),
   561 => (x"a6",x"c8",x"87",x"c8"),
   562 => (x"c0",x"78",x"c0",x"48"),
   563 => (x"a6",x"c8",x"87",x"c5"),
   564 => (x"c8",x"78",x"c1",x"48"),
   565 => (x"9c",x"74",x"4c",x"66"),
   566 => (x"87",x"e0",x"c0",x"05"),
   567 => (x"c2",x"49",x"66",x"c4"),
   568 => (x"c4",x"c9",x"c2",x"89"),
   569 => (x"c2",x"91",x"4a",x"bf"),
   570 => (x"4a",x"bf",x"dd",x"cd"),
   571 => (x"48",x"f8",x"c0",x"c2"),
   572 => (x"c2",x"78",x"a1",x"72"),
   573 => (x"c0",x"48",x"c0",x"c1"),
   574 => (x"87",x"e1",x"f9",x"78"),
   575 => (x"8e",x"f4",x"48",x"c0"),
   576 => (x"00",x"87",x"d9",x"ee"),
   577 => (x"ff",x"00",x"00",x"00"),
   578 => (x"13",x"ff",x"ff",x"ff"),
   579 => (x"1c",x"00",x"00",x"09"),
   580 => (x"46",x"00",x"00",x"09"),
   581 => (x"32",x"33",x"54",x"41"),
   582 => (x"00",x"20",x"20",x"20"),
   583 => (x"31",x"54",x"41",x"46"),
   584 => (x"20",x"20",x"20",x"36"),
   585 => (x"d4",x"ff",x"1e",x"00"),
   586 => (x"78",x"ff",x"c3",x"48"),
   587 => (x"4f",x"26",x"48",x"68"),
   588 => (x"48",x"d4",x"ff",x"1e"),
   589 => (x"ff",x"78",x"ff",x"c3"),
   590 => (x"e1",x"c0",x"48",x"d0"),
   591 => (x"48",x"d4",x"ff",x"78"),
   592 => (x"cd",x"c2",x"78",x"d4"),
   593 => (x"d4",x"ff",x"48",x"f5"),
   594 => (x"4f",x"26",x"50",x"bf"),
   595 => (x"48",x"d0",x"ff",x"1e"),
   596 => (x"26",x"78",x"e0",x"c0"),
   597 => (x"cc",x"ff",x"1e",x"4f"),
   598 => (x"99",x"49",x"70",x"87"),
   599 => (x"c0",x"87",x"c6",x"02"),
   600 => (x"f1",x"05",x"a9",x"fb"),
   601 => (x"26",x"48",x"71",x"87"),
   602 => (x"5b",x"5e",x"0e",x"4f"),
   603 => (x"4b",x"71",x"0e",x"5c"),
   604 => (x"f0",x"fe",x"4c",x"c0"),
   605 => (x"99",x"49",x"70",x"87"),
   606 => (x"87",x"f9",x"c0",x"02"),
   607 => (x"02",x"a9",x"ec",x"c0"),
   608 => (x"c0",x"87",x"f2",x"c0"),
   609 => (x"c0",x"02",x"a9",x"fb"),
   610 => (x"66",x"cc",x"87",x"eb"),
   611 => (x"c7",x"03",x"ac",x"b7"),
   612 => (x"02",x"66",x"d0",x"87"),
   613 => (x"53",x"71",x"87",x"c2"),
   614 => (x"c2",x"02",x"99",x"71"),
   615 => (x"fe",x"84",x"c1",x"87"),
   616 => (x"49",x"70",x"87",x"c3"),
   617 => (x"87",x"cd",x"02",x"99"),
   618 => (x"02",x"a9",x"ec",x"c0"),
   619 => (x"fb",x"c0",x"87",x"c7"),
   620 => (x"d5",x"ff",x"05",x"a9"),
   621 => (x"02",x"66",x"d0",x"87"),
   622 => (x"97",x"c0",x"87",x"c3"),
   623 => (x"a9",x"ec",x"c0",x"7b"),
   624 => (x"74",x"87",x"c4",x"05"),
   625 => (x"74",x"87",x"c5",x"4a"),
   626 => (x"8a",x"0a",x"c0",x"4a"),
   627 => (x"87",x"c2",x"48",x"72"),
   628 => (x"4c",x"26",x"4d",x"26"),
   629 => (x"4f",x"26",x"4b",x"26"),
   630 => (x"87",x"c9",x"fd",x"1e"),
   631 => (x"c0",x"4a",x"49",x"70"),
   632 => (x"c9",x"04",x"aa",x"f0"),
   633 => (x"aa",x"f9",x"c0",x"87"),
   634 => (x"c0",x"87",x"c3",x"01"),
   635 => (x"c1",x"c1",x"8a",x"f0"),
   636 => (x"87",x"c9",x"04",x"aa"),
   637 => (x"01",x"aa",x"da",x"c1"),
   638 => (x"f7",x"c0",x"87",x"c3"),
   639 => (x"26",x"48",x"72",x"8a"),
   640 => (x"5b",x"5e",x"0e",x"4f"),
   641 => (x"4a",x"71",x"0e",x"5c"),
   642 => (x"72",x"4b",x"d4",x"ff"),
   643 => (x"87",x"e7",x"c0",x"49"),
   644 => (x"02",x"9c",x"4c",x"70"),
   645 => (x"8c",x"c1",x"87",x"c2"),
   646 => (x"c5",x"48",x"d0",x"ff"),
   647 => (x"7b",x"d5",x"c1",x"78"),
   648 => (x"31",x"c6",x"49",x"74"),
   649 => (x"97",x"f7",x"d2",x"c1"),
   650 => (x"71",x"48",x"4a",x"bf"),
   651 => (x"ff",x"7b",x"70",x"b0"),
   652 => (x"78",x"c4",x"48",x"d0"),
   653 => (x"0e",x"87",x"db",x"fe"),
   654 => (x"5d",x"5c",x"5b",x"5e"),
   655 => (x"71",x"86",x"f8",x"0e"),
   656 => (x"fb",x"7e",x"c0",x"4c"),
   657 => (x"4b",x"c0",x"87",x"ea"),
   658 => (x"97",x"e4",x"eb",x"c0"),
   659 => (x"a9",x"c0",x"49",x"bf"),
   660 => (x"fb",x"87",x"cf",x"04"),
   661 => (x"83",x"c1",x"87",x"ff"),
   662 => (x"97",x"e4",x"eb",x"c0"),
   663 => (x"06",x"ab",x"49",x"bf"),
   664 => (x"eb",x"c0",x"87",x"f1"),
   665 => (x"02",x"bf",x"97",x"e4"),
   666 => (x"f8",x"fa",x"87",x"cf"),
   667 => (x"99",x"49",x"70",x"87"),
   668 => (x"c0",x"87",x"c6",x"02"),
   669 => (x"f1",x"05",x"a9",x"ec"),
   670 => (x"fa",x"4b",x"c0",x"87"),
   671 => (x"4d",x"70",x"87",x"e7"),
   672 => (x"c8",x"87",x"e2",x"fa"),
   673 => (x"dc",x"fa",x"58",x"a6"),
   674 => (x"c1",x"4a",x"70",x"87"),
   675 => (x"49",x"a4",x"c8",x"83"),
   676 => (x"ad",x"49",x"69",x"97"),
   677 => (x"c0",x"87",x"c7",x"02"),
   678 => (x"c0",x"05",x"ad",x"ff"),
   679 => (x"a4",x"c9",x"87",x"e7"),
   680 => (x"49",x"69",x"97",x"49"),
   681 => (x"02",x"a9",x"66",x"c4"),
   682 => (x"c0",x"48",x"87",x"c7"),
   683 => (x"d4",x"05",x"a8",x"ff"),
   684 => (x"49",x"a4",x"ca",x"87"),
   685 => (x"aa",x"49",x"69",x"97"),
   686 => (x"c0",x"87",x"c6",x"02"),
   687 => (x"c4",x"05",x"aa",x"ff"),
   688 => (x"d0",x"7e",x"c1",x"87"),
   689 => (x"ad",x"ec",x"c0",x"87"),
   690 => (x"c0",x"87",x"c6",x"02"),
   691 => (x"c4",x"05",x"ad",x"fb"),
   692 => (x"c1",x"4b",x"c0",x"87"),
   693 => (x"fe",x"02",x"6e",x"7e"),
   694 => (x"ef",x"f9",x"87",x"e1"),
   695 => (x"f8",x"48",x"73",x"87"),
   696 => (x"87",x"ec",x"fb",x"8e"),
   697 => (x"5b",x"5e",x"0e",x"00"),
   698 => (x"f8",x"0e",x"5d",x"5c"),
   699 => (x"ff",x"4d",x"71",x"86"),
   700 => (x"1e",x"75",x"4b",x"d4"),
   701 => (x"49",x"fa",x"cd",x"c2"),
   702 => (x"c4",x"87",x"db",x"e8"),
   703 => (x"02",x"98",x"70",x"86"),
   704 => (x"c4",x"87",x"cc",x"c4"),
   705 => (x"d2",x"c1",x"48",x"a6"),
   706 => (x"75",x"78",x"bf",x"f9"),
   707 => (x"87",x"f1",x"fb",x"49"),
   708 => (x"c5",x"48",x"d0",x"ff"),
   709 => (x"7b",x"d6",x"c1",x"78"),
   710 => (x"a2",x"75",x"4a",x"c0"),
   711 => (x"c1",x"7b",x"11",x"49"),
   712 => (x"aa",x"b7",x"cb",x"82"),
   713 => (x"cc",x"87",x"f3",x"04"),
   714 => (x"7b",x"ff",x"c3",x"4a"),
   715 => (x"e0",x"c0",x"82",x"c1"),
   716 => (x"f4",x"04",x"aa",x"b7"),
   717 => (x"48",x"d0",x"ff",x"87"),
   718 => (x"ff",x"c3",x"78",x"c4"),
   719 => (x"c1",x"78",x"c5",x"7b"),
   720 => (x"7b",x"c1",x"7b",x"d3"),
   721 => (x"48",x"66",x"78",x"c4"),
   722 => (x"06",x"a8",x"b7",x"c0"),
   723 => (x"c2",x"87",x"f0",x"c2"),
   724 => (x"4c",x"bf",x"c2",x"ce"),
   725 => (x"74",x"48",x"66",x"c4"),
   726 => (x"58",x"a6",x"c8",x"88"),
   727 => (x"c1",x"02",x"9c",x"74"),
   728 => (x"c1",x"c2",x"87",x"f9"),
   729 => (x"c0",x"c8",x"7e",x"c4"),
   730 => (x"b7",x"c0",x"8c",x"4d"),
   731 => (x"87",x"c6",x"03",x"ac"),
   732 => (x"4d",x"a4",x"c0",x"c8"),
   733 => (x"cd",x"c2",x"4c",x"c0"),
   734 => (x"49",x"bf",x"97",x"f5"),
   735 => (x"d1",x"02",x"99",x"d0"),
   736 => (x"c2",x"1e",x"c0",x"87"),
   737 => (x"ea",x"49",x"fa",x"cd"),
   738 => (x"86",x"c4",x"87",x"ff"),
   739 => (x"c0",x"4a",x"49",x"70"),
   740 => (x"c1",x"c2",x"87",x"ee"),
   741 => (x"cd",x"c2",x"1e",x"c4"),
   742 => (x"ec",x"ea",x"49",x"fa"),
   743 => (x"70",x"86",x"c4",x"87"),
   744 => (x"d0",x"ff",x"4a",x"49"),
   745 => (x"78",x"c5",x"c8",x"48"),
   746 => (x"6e",x"7b",x"d4",x"c1"),
   747 => (x"6e",x"7b",x"bf",x"97"),
   748 => (x"70",x"80",x"c1",x"48"),
   749 => (x"05",x"8d",x"c1",x"7e"),
   750 => (x"ff",x"87",x"f0",x"ff"),
   751 => (x"78",x"c4",x"48",x"d0"),
   752 => (x"c5",x"05",x"9a",x"72"),
   753 => (x"c1",x"48",x"c0",x"87"),
   754 => (x"1e",x"c1",x"87",x"c7"),
   755 => (x"49",x"fa",x"cd",x"c2"),
   756 => (x"c4",x"87",x"dc",x"e8"),
   757 => (x"05",x"9c",x"74",x"86"),
   758 => (x"c4",x"87",x"c7",x"fe"),
   759 => (x"b7",x"c0",x"48",x"66"),
   760 => (x"87",x"d1",x"06",x"a8"),
   761 => (x"48",x"fa",x"cd",x"c2"),
   762 => (x"80",x"d0",x"78",x"c0"),
   763 => (x"80",x"f4",x"78",x"c0"),
   764 => (x"bf",x"c6",x"ce",x"c2"),
   765 => (x"48",x"66",x"c4",x"78"),
   766 => (x"01",x"a8",x"b7",x"c0"),
   767 => (x"ff",x"87",x"d0",x"fd"),
   768 => (x"78",x"c5",x"48",x"d0"),
   769 => (x"c0",x"7b",x"d3",x"c1"),
   770 => (x"c1",x"78",x"c4",x"7b"),
   771 => (x"c0",x"87",x"c2",x"48"),
   772 => (x"26",x"8e",x"f8",x"48"),
   773 => (x"26",x"4c",x"26",x"4d"),
   774 => (x"0e",x"4f",x"26",x"4b"),
   775 => (x"5d",x"5c",x"5b",x"5e"),
   776 => (x"4b",x"71",x"1e",x"0e"),
   777 => (x"ab",x"4d",x"4c",x"c0"),
   778 => (x"87",x"e8",x"c0",x"04"),
   779 => (x"1e",x"f7",x"e8",x"c0"),
   780 => (x"c4",x"02",x"9d",x"75"),
   781 => (x"c2",x"4a",x"c0",x"87"),
   782 => (x"72",x"4a",x"c1",x"87"),
   783 => (x"87",x"ee",x"eb",x"49"),
   784 => (x"7e",x"70",x"86",x"c4"),
   785 => (x"05",x"6e",x"84",x"c1"),
   786 => (x"4c",x"73",x"87",x"c2"),
   787 => (x"ac",x"73",x"85",x"c1"),
   788 => (x"87",x"d8",x"ff",x"06"),
   789 => (x"fe",x"26",x"48",x"6e"),
   790 => (x"71",x"1e",x"87",x"f9"),
   791 => (x"05",x"66",x"c4",x"4a"),
   792 => (x"49",x"72",x"87",x"c5"),
   793 => (x"26",x"87",x"fe",x"f9"),
   794 => (x"5b",x"5e",x"0e",x"4f"),
   795 => (x"1e",x"0e",x"5d",x"5c"),
   796 => (x"de",x"49",x"4c",x"71"),
   797 => (x"e2",x"ce",x"c2",x"91"),
   798 => (x"97",x"85",x"71",x"4d"),
   799 => (x"dd",x"c1",x"02",x"6d"),
   800 => (x"ce",x"ce",x"c2",x"87"),
   801 => (x"82",x"74",x"4a",x"bf"),
   802 => (x"ce",x"fe",x"49",x"72"),
   803 => (x"48",x"7e",x"70",x"87"),
   804 => (x"f2",x"c0",x"02",x"98"),
   805 => (x"d6",x"ce",x"c2",x"87"),
   806 => (x"cb",x"4a",x"70",x"4b"),
   807 => (x"c6",x"d0",x"ff",x"49"),
   808 => (x"cb",x"4b",x"74",x"87"),
   809 => (x"cb",x"d3",x"c1",x"93"),
   810 => (x"c0",x"83",x"c4",x"83"),
   811 => (x"74",x"7b",x"e2",x"f3"),
   812 => (x"df",x"fe",x"c0",x"49"),
   813 => (x"c1",x"7b",x"75",x"87"),
   814 => (x"bf",x"97",x"f8",x"d2"),
   815 => (x"ce",x"c2",x"1e",x"49"),
   816 => (x"d5",x"fe",x"49",x"d6"),
   817 => (x"74",x"86",x"c4",x"87"),
   818 => (x"c7",x"fe",x"c0",x"49"),
   819 => (x"c0",x"49",x"c0",x"87"),
   820 => (x"c2",x"87",x"e6",x"ff"),
   821 => (x"c0",x"48",x"f6",x"cd"),
   822 => (x"de",x"49",x"c1",x"78"),
   823 => (x"fc",x"26",x"87",x"dc"),
   824 => (x"6f",x"4c",x"87",x"f1"),
   825 => (x"6e",x"69",x"64",x"61"),
   826 => (x"2e",x"2e",x"2e",x"67"),
   827 => (x"5b",x"5e",x"0e",x"00"),
   828 => (x"4b",x"71",x"0e",x"5c"),
   829 => (x"ce",x"ce",x"c2",x"4a"),
   830 => (x"49",x"72",x"82",x"bf"),
   831 => (x"70",x"87",x"dc",x"fc"),
   832 => (x"c4",x"02",x"9c",x"4c"),
   833 => (x"ed",x"e7",x"49",x"87"),
   834 => (x"ce",x"ce",x"c2",x"87"),
   835 => (x"c1",x"78",x"c0",x"48"),
   836 => (x"87",x"e6",x"dd",x"49"),
   837 => (x"0e",x"87",x"fe",x"fb"),
   838 => (x"5d",x"5c",x"5b",x"5e"),
   839 => (x"c2",x"86",x"f4",x"0e"),
   840 => (x"c0",x"4d",x"c4",x"c1"),
   841 => (x"48",x"a6",x"c4",x"4c"),
   842 => (x"ce",x"c2",x"78",x"c0"),
   843 => (x"c0",x"49",x"bf",x"ce"),
   844 => (x"c1",x"c1",x"06",x"a9"),
   845 => (x"c4",x"c1",x"c2",x"87"),
   846 => (x"c0",x"02",x"98",x"48"),
   847 => (x"e8",x"c0",x"87",x"f8"),
   848 => (x"66",x"c8",x"1e",x"f7"),
   849 => (x"c4",x"87",x"c7",x"02"),
   850 => (x"78",x"c0",x"48",x"a6"),
   851 => (x"a6",x"c4",x"87",x"c5"),
   852 => (x"c4",x"78",x"c1",x"48"),
   853 => (x"d5",x"e7",x"49",x"66"),
   854 => (x"70",x"86",x"c4",x"87"),
   855 => (x"c4",x"84",x"c1",x"4d"),
   856 => (x"80",x"c1",x"48",x"66"),
   857 => (x"c2",x"58",x"a6",x"c8"),
   858 => (x"49",x"bf",x"ce",x"ce"),
   859 => (x"87",x"c6",x"03",x"ac"),
   860 => (x"ff",x"05",x"9d",x"75"),
   861 => (x"4c",x"c0",x"87",x"c8"),
   862 => (x"c3",x"02",x"9d",x"75"),
   863 => (x"e8",x"c0",x"87",x"e0"),
   864 => (x"66",x"c8",x"1e",x"f7"),
   865 => (x"cc",x"87",x"c7",x"02"),
   866 => (x"78",x"c0",x"48",x"a6"),
   867 => (x"a6",x"cc",x"87",x"c5"),
   868 => (x"cc",x"78",x"c1",x"48"),
   869 => (x"d5",x"e6",x"49",x"66"),
   870 => (x"70",x"86",x"c4",x"87"),
   871 => (x"02",x"98",x"48",x"7e"),
   872 => (x"49",x"87",x"e8",x"c2"),
   873 => (x"69",x"97",x"81",x"cb"),
   874 => (x"02",x"99",x"d0",x"49"),
   875 => (x"c0",x"87",x"d6",x"c1"),
   876 => (x"74",x"4a",x"ed",x"f3"),
   877 => (x"c1",x"91",x"cb",x"49"),
   878 => (x"72",x"81",x"cb",x"d3"),
   879 => (x"c3",x"81",x"c8",x"79"),
   880 => (x"49",x"74",x"51",x"ff"),
   881 => (x"ce",x"c2",x"91",x"de"),
   882 => (x"85",x"71",x"4d",x"e2"),
   883 => (x"7d",x"97",x"c1",x"c2"),
   884 => (x"c0",x"49",x"a5",x"c1"),
   885 => (x"c9",x"c2",x"51",x"e0"),
   886 => (x"02",x"bf",x"97",x"d4"),
   887 => (x"84",x"c1",x"87",x"d2"),
   888 => (x"c2",x"4b",x"a5",x"c2"),
   889 => (x"db",x"4a",x"d4",x"c9"),
   890 => (x"fa",x"ca",x"ff",x"49"),
   891 => (x"87",x"db",x"c1",x"87"),
   892 => (x"c0",x"49",x"a5",x"cd"),
   893 => (x"c2",x"84",x"c1",x"51"),
   894 => (x"4a",x"6e",x"4b",x"a5"),
   895 => (x"ca",x"ff",x"49",x"cb"),
   896 => (x"c6",x"c1",x"87",x"e5"),
   897 => (x"e9",x"f1",x"c0",x"87"),
   898 => (x"cb",x"49",x"74",x"4a"),
   899 => (x"cb",x"d3",x"c1",x"91"),
   900 => (x"c2",x"79",x"72",x"81"),
   901 => (x"bf",x"97",x"d4",x"c9"),
   902 => (x"74",x"87",x"d8",x"02"),
   903 => (x"c1",x"91",x"de",x"49"),
   904 => (x"e2",x"ce",x"c2",x"84"),
   905 => (x"c2",x"83",x"71",x"4b"),
   906 => (x"dd",x"4a",x"d4",x"c9"),
   907 => (x"f6",x"c9",x"ff",x"49"),
   908 => (x"74",x"87",x"d8",x"87"),
   909 => (x"c2",x"93",x"de",x"4b"),
   910 => (x"cb",x"83",x"e2",x"ce"),
   911 => (x"51",x"c0",x"49",x"a3"),
   912 => (x"6e",x"73",x"84",x"c1"),
   913 => (x"ff",x"49",x"cb",x"4a"),
   914 => (x"c4",x"87",x"dc",x"c9"),
   915 => (x"80",x"c1",x"48",x"66"),
   916 => (x"c7",x"58",x"a6",x"c8"),
   917 => (x"c5",x"c0",x"03",x"ac"),
   918 => (x"fc",x"05",x"6e",x"87"),
   919 => (x"48",x"74",x"87",x"e0"),
   920 => (x"ee",x"f6",x"8e",x"f4"),
   921 => (x"1e",x"73",x"1e",x"87"),
   922 => (x"cb",x"49",x"4b",x"71"),
   923 => (x"cb",x"d3",x"c1",x"91"),
   924 => (x"4a",x"a1",x"c8",x"81"),
   925 => (x"48",x"f7",x"d2",x"c1"),
   926 => (x"a1",x"c9",x"50",x"12"),
   927 => (x"e4",x"eb",x"c0",x"4a"),
   928 => (x"ca",x"50",x"12",x"48"),
   929 => (x"f8",x"d2",x"c1",x"81"),
   930 => (x"c1",x"50",x"11",x"48"),
   931 => (x"bf",x"97",x"f8",x"d2"),
   932 => (x"49",x"c0",x"1e",x"49"),
   933 => (x"c2",x"87",x"c3",x"f7"),
   934 => (x"de",x"48",x"f6",x"cd"),
   935 => (x"d7",x"49",x"c1",x"78"),
   936 => (x"f5",x"26",x"87",x"d8"),
   937 => (x"71",x"1e",x"87",x"f1"),
   938 => (x"91",x"cb",x"49",x"4a"),
   939 => (x"81",x"cb",x"d3",x"c1"),
   940 => (x"48",x"11",x"81",x"c8"),
   941 => (x"58",x"fa",x"cd",x"c2"),
   942 => (x"48",x"ce",x"ce",x"c2"),
   943 => (x"49",x"c1",x"78",x"c0"),
   944 => (x"26",x"87",x"f7",x"d6"),
   945 => (x"49",x"c0",x"1e",x"4f"),
   946 => (x"87",x"ed",x"f7",x"c0"),
   947 => (x"71",x"1e",x"4f",x"26"),
   948 => (x"87",x"d2",x"02",x"99"),
   949 => (x"48",x"e0",x"d4",x"c1"),
   950 => (x"80",x"f7",x"50",x"c0"),
   951 => (x"40",x"e6",x"fa",x"c0"),
   952 => (x"78",x"c4",x"d3",x"c1"),
   953 => (x"d4",x"c1",x"87",x"ce"),
   954 => (x"d2",x"c1",x"48",x"dc"),
   955 => (x"80",x"fc",x"78",x"fd"),
   956 => (x"78",x"c5",x"fb",x"c0"),
   957 => (x"5e",x"0e",x"4f",x"26"),
   958 => (x"0e",x"5d",x"5c",x"5b"),
   959 => (x"4d",x"71",x"86",x"f4"),
   960 => (x"c1",x"91",x"cb",x"49"),
   961 => (x"c8",x"81",x"cb",x"d3"),
   962 => (x"a1",x"ca",x"4a",x"a1"),
   963 => (x"48",x"a6",x"c4",x"7e"),
   964 => (x"bf",x"fe",x"d1",x"c2"),
   965 => (x"bf",x"97",x"6e",x"78"),
   966 => (x"48",x"66",x"c4",x"4b"),
   967 => (x"4b",x"70",x"28",x"73"),
   968 => (x"cc",x"48",x"12",x"4c"),
   969 => (x"9c",x"70",x"58",x"a6"),
   970 => (x"81",x"c9",x"84",x"c1"),
   971 => (x"b7",x"49",x"69",x"97"),
   972 => (x"87",x"c2",x"04",x"ac"),
   973 => (x"97",x"6e",x"4c",x"c0"),
   974 => (x"66",x"c8",x"4a",x"bf"),
   975 => (x"ff",x"31",x"72",x"49"),
   976 => (x"99",x"66",x"c4",x"b9"),
   977 => (x"30",x"72",x"48",x"74"),
   978 => (x"71",x"48",x"4a",x"70"),
   979 => (x"c2",x"d2",x"c2",x"b0"),
   980 => (x"ff",x"e1",x"c0",x"58"),
   981 => (x"d4",x"49",x"c0",x"87"),
   982 => (x"49",x"75",x"87",x"e0"),
   983 => (x"87",x"f4",x"f3",x"c0"),
   984 => (x"ee",x"f2",x"8e",x"f4"),
   985 => (x"1e",x"73",x"1e",x"87"),
   986 => (x"fe",x"49",x"4b",x"71"),
   987 => (x"49",x"73",x"87",x"c8"),
   988 => (x"f2",x"87",x"c3",x"fe"),
   989 => (x"73",x"1e",x"87",x"e1"),
   990 => (x"c6",x"4b",x"71",x"1e"),
   991 => (x"db",x"02",x"4a",x"a3"),
   992 => (x"02",x"8a",x"c1",x"87"),
   993 => (x"02",x"8a",x"87",x"d6"),
   994 => (x"8a",x"87",x"da",x"c1"),
   995 => (x"87",x"fc",x"c0",x"02"),
   996 => (x"e1",x"c0",x"02",x"8a"),
   997 => (x"cb",x"02",x"8a",x"87"),
   998 => (x"87",x"db",x"c1",x"87"),
   999 => (x"c5",x"fc",x"49",x"c7"),
  1000 => (x"87",x"de",x"c1",x"87"),
  1001 => (x"bf",x"ce",x"ce",x"c2"),
  1002 => (x"87",x"cb",x"c1",x"02"),
  1003 => (x"c2",x"88",x"c1",x"48"),
  1004 => (x"c1",x"58",x"d2",x"ce"),
  1005 => (x"ce",x"c2",x"87",x"c1"),
  1006 => (x"c0",x"02",x"bf",x"d2"),
  1007 => (x"ce",x"c2",x"87",x"f9"),
  1008 => (x"c1",x"48",x"bf",x"ce"),
  1009 => (x"d2",x"ce",x"c2",x"80"),
  1010 => (x"87",x"eb",x"c0",x"58"),
  1011 => (x"bf",x"ce",x"ce",x"c2"),
  1012 => (x"c2",x"89",x"c6",x"49"),
  1013 => (x"c0",x"59",x"d2",x"ce"),
  1014 => (x"da",x"03",x"a9",x"b7"),
  1015 => (x"ce",x"ce",x"c2",x"87"),
  1016 => (x"d2",x"78",x"c0",x"48"),
  1017 => (x"d2",x"ce",x"c2",x"87"),
  1018 => (x"87",x"cb",x"02",x"bf"),
  1019 => (x"bf",x"ce",x"ce",x"c2"),
  1020 => (x"c2",x"80",x"c6",x"48"),
  1021 => (x"c0",x"58",x"d2",x"ce"),
  1022 => (x"87",x"fe",x"d1",x"49"),
  1023 => (x"f1",x"c0",x"49",x"73"),
  1024 => (x"d2",x"f0",x"87",x"d2"),
  1025 => (x"5b",x"5e",x"0e",x"87"),
  1026 => (x"ff",x"0e",x"5d",x"5c"),
  1027 => (x"a6",x"dc",x"86",x"d0"),
  1028 => (x"48",x"a6",x"c8",x"59"),
  1029 => (x"80",x"c4",x"78",x"c0"),
  1030 => (x"78",x"66",x"c4",x"c1"),
  1031 => (x"78",x"c1",x"80",x"c4"),
  1032 => (x"78",x"c1",x"80",x"c4"),
  1033 => (x"48",x"d2",x"ce",x"c2"),
  1034 => (x"cd",x"c2",x"78",x"c1"),
  1035 => (x"de",x"48",x"bf",x"f6"),
  1036 => (x"87",x"cb",x"05",x"a8"),
  1037 => (x"70",x"87",x"e0",x"f3"),
  1038 => (x"59",x"a6",x"cc",x"49"),
  1039 => (x"e3",x"87",x"fa",x"cf"),
  1040 => (x"d0",x"e4",x"87",x"ee"),
  1041 => (x"87",x"dd",x"e3",x"87"),
  1042 => (x"fb",x"c0",x"4c",x"70"),
  1043 => (x"fb",x"c1",x"02",x"ac"),
  1044 => (x"05",x"66",x"d8",x"87"),
  1045 => (x"c1",x"87",x"ed",x"c1"),
  1046 => (x"c4",x"4a",x"66",x"c0"),
  1047 => (x"72",x"7e",x"6a",x"82"),
  1048 => (x"ee",x"d1",x"c1",x"1e"),
  1049 => (x"49",x"66",x"c4",x"48"),
  1050 => (x"20",x"4a",x"a1",x"c8"),
  1051 => (x"05",x"aa",x"71",x"41"),
  1052 => (x"51",x"10",x"87",x"f9"),
  1053 => (x"c0",x"c1",x"4a",x"26"),
  1054 => (x"f9",x"c0",x"48",x"66"),
  1055 => (x"49",x"6a",x"78",x"e5"),
  1056 => (x"51",x"74",x"81",x"c7"),
  1057 => (x"49",x"66",x"c0",x"c1"),
  1058 => (x"51",x"c1",x"81",x"c8"),
  1059 => (x"49",x"66",x"c0",x"c1"),
  1060 => (x"51",x"c0",x"81",x"c9"),
  1061 => (x"49",x"66",x"c0",x"c1"),
  1062 => (x"51",x"c0",x"81",x"ca"),
  1063 => (x"1e",x"d8",x"1e",x"c1"),
  1064 => (x"81",x"c8",x"49",x"6a"),
  1065 => (x"c8",x"87",x"c2",x"e3"),
  1066 => (x"66",x"c4",x"c1",x"86"),
  1067 => (x"01",x"a8",x"c0",x"48"),
  1068 => (x"a6",x"c8",x"87",x"c7"),
  1069 => (x"ce",x"78",x"c1",x"48"),
  1070 => (x"66",x"c4",x"c1",x"87"),
  1071 => (x"d0",x"88",x"c1",x"48"),
  1072 => (x"87",x"c3",x"58",x"a6"),
  1073 => (x"d0",x"87",x"ce",x"e2"),
  1074 => (x"78",x"c2",x"48",x"a6"),
  1075 => (x"cd",x"02",x"9c",x"74"),
  1076 => (x"66",x"c8",x"87",x"e3"),
  1077 => (x"66",x"c8",x"c1",x"48"),
  1078 => (x"d8",x"cd",x"03",x"a8"),
  1079 => (x"48",x"a6",x"dc",x"87"),
  1080 => (x"80",x"e8",x"78",x"c0"),
  1081 => (x"fc",x"e0",x"78",x"c0"),
  1082 => (x"c1",x"4c",x"70",x"87"),
  1083 => (x"c2",x"05",x"ac",x"d0"),
  1084 => (x"66",x"c4",x"87",x"d8"),
  1085 => (x"87",x"e0",x"e3",x"7e"),
  1086 => (x"a6",x"c8",x"49",x"70"),
  1087 => (x"87",x"e5",x"e0",x"59"),
  1088 => (x"ec",x"c0",x"4c",x"70"),
  1089 => (x"ec",x"c1",x"05",x"ac"),
  1090 => (x"49",x"66",x"c8",x"87"),
  1091 => (x"c0",x"c1",x"91",x"cb"),
  1092 => (x"a1",x"c4",x"81",x"66"),
  1093 => (x"c8",x"4d",x"6a",x"4a"),
  1094 => (x"66",x"c4",x"4a",x"a1"),
  1095 => (x"e6",x"fa",x"c0",x"52"),
  1096 => (x"87",x"c1",x"e0",x"79"),
  1097 => (x"02",x"9c",x"4c",x"70"),
  1098 => (x"fb",x"c0",x"87",x"d9"),
  1099 => (x"87",x"d3",x"02",x"ac"),
  1100 => (x"df",x"ff",x"55",x"74"),
  1101 => (x"4c",x"70",x"87",x"ef"),
  1102 => (x"87",x"c7",x"02",x"9c"),
  1103 => (x"05",x"ac",x"fb",x"c0"),
  1104 => (x"c0",x"87",x"ed",x"ff"),
  1105 => (x"c1",x"c2",x"55",x"e0"),
  1106 => (x"7d",x"97",x"c0",x"55"),
  1107 => (x"6e",x"49",x"66",x"d8"),
  1108 => (x"87",x"db",x"05",x"a9"),
  1109 => (x"cc",x"48",x"66",x"c8"),
  1110 => (x"ca",x"04",x"a8",x"66"),
  1111 => (x"48",x"66",x"c8",x"87"),
  1112 => (x"a6",x"cc",x"80",x"c1"),
  1113 => (x"cc",x"87",x"c8",x"58"),
  1114 => (x"88",x"c1",x"48",x"66"),
  1115 => (x"ff",x"58",x"a6",x"d0"),
  1116 => (x"70",x"87",x"f2",x"de"),
  1117 => (x"ac",x"d0",x"c1",x"4c"),
  1118 => (x"d4",x"87",x"c8",x"05"),
  1119 => (x"80",x"c1",x"48",x"66"),
  1120 => (x"c1",x"58",x"a6",x"d8"),
  1121 => (x"fd",x"02",x"ac",x"d0"),
  1122 => (x"e0",x"c0",x"87",x"e8"),
  1123 => (x"66",x"d8",x"48",x"a6"),
  1124 => (x"48",x"66",x"c4",x"78"),
  1125 => (x"a8",x"66",x"e0",x"c0"),
  1126 => (x"87",x"eb",x"c9",x"05"),
  1127 => (x"48",x"a6",x"e4",x"c0"),
  1128 => (x"48",x"74",x"78",x"c0"),
  1129 => (x"70",x"88",x"fb",x"c0"),
  1130 => (x"02",x"98",x"48",x"7e"),
  1131 => (x"48",x"87",x"ed",x"c9"),
  1132 => (x"7e",x"70",x"88",x"cb"),
  1133 => (x"c1",x"02",x"98",x"48"),
  1134 => (x"c9",x"48",x"87",x"cd"),
  1135 => (x"48",x"7e",x"70",x"88"),
  1136 => (x"c1",x"c4",x"02",x"98"),
  1137 => (x"88",x"c4",x"48",x"87"),
  1138 => (x"98",x"48",x"7e",x"70"),
  1139 => (x"48",x"87",x"ce",x"02"),
  1140 => (x"7e",x"70",x"88",x"c1"),
  1141 => (x"c3",x"02",x"98",x"48"),
  1142 => (x"e1",x"c8",x"87",x"ec"),
  1143 => (x"48",x"a6",x"dc",x"87"),
  1144 => (x"ff",x"78",x"f0",x"c0"),
  1145 => (x"70",x"87",x"fe",x"dc"),
  1146 => (x"ac",x"ec",x"c0",x"4c"),
  1147 => (x"87",x"c4",x"c0",x"02"),
  1148 => (x"5c",x"a6",x"e0",x"c0"),
  1149 => (x"02",x"ac",x"ec",x"c0"),
  1150 => (x"dc",x"ff",x"87",x"cd"),
  1151 => (x"4c",x"70",x"87",x"e7"),
  1152 => (x"05",x"ac",x"ec",x"c0"),
  1153 => (x"c0",x"87",x"f3",x"ff"),
  1154 => (x"c0",x"02",x"ac",x"ec"),
  1155 => (x"dc",x"ff",x"87",x"c4"),
  1156 => (x"1e",x"c0",x"87",x"d3"),
  1157 => (x"66",x"d0",x"1e",x"ca"),
  1158 => (x"c1",x"91",x"cb",x"49"),
  1159 => (x"71",x"48",x"66",x"c8"),
  1160 => (x"58",x"a6",x"cc",x"80"),
  1161 => (x"c4",x"48",x"66",x"c8"),
  1162 => (x"58",x"a6",x"d0",x"80"),
  1163 => (x"49",x"bf",x"66",x"cc"),
  1164 => (x"87",x"f5",x"dc",x"ff"),
  1165 => (x"1e",x"de",x"1e",x"c1"),
  1166 => (x"49",x"bf",x"66",x"d4"),
  1167 => (x"87",x"e9",x"dc",x"ff"),
  1168 => (x"49",x"70",x"86",x"d0"),
  1169 => (x"c0",x"89",x"09",x"c0"),
  1170 => (x"c0",x"59",x"a6",x"ec"),
  1171 => (x"c0",x"48",x"66",x"e8"),
  1172 => (x"ee",x"c0",x"06",x"a8"),
  1173 => (x"66",x"e8",x"c0",x"87"),
  1174 => (x"03",x"a8",x"dd",x"48"),
  1175 => (x"c4",x"87",x"e4",x"c0"),
  1176 => (x"c0",x"49",x"bf",x"66"),
  1177 => (x"c0",x"81",x"66",x"e8"),
  1178 => (x"e8",x"c0",x"51",x"e0"),
  1179 => (x"81",x"c1",x"49",x"66"),
  1180 => (x"81",x"bf",x"66",x"c4"),
  1181 => (x"c0",x"51",x"c1",x"c2"),
  1182 => (x"c2",x"49",x"66",x"e8"),
  1183 => (x"bf",x"66",x"c4",x"81"),
  1184 => (x"6e",x"51",x"c0",x"81"),
  1185 => (x"e5",x"f9",x"c0",x"48"),
  1186 => (x"c8",x"49",x"6e",x"78"),
  1187 => (x"51",x"66",x"d0",x"81"),
  1188 => (x"81",x"c9",x"49",x"6e"),
  1189 => (x"6e",x"51",x"66",x"d4"),
  1190 => (x"dc",x"81",x"ca",x"49"),
  1191 => (x"66",x"d0",x"51",x"66"),
  1192 => (x"d4",x"80",x"c1",x"48"),
  1193 => (x"66",x"c8",x"58",x"a6"),
  1194 => (x"a8",x"66",x"cc",x"48"),
  1195 => (x"87",x"cb",x"c0",x"04"),
  1196 => (x"c1",x"48",x"66",x"c8"),
  1197 => (x"58",x"a6",x"cc",x"80"),
  1198 => (x"cc",x"87",x"e1",x"c5"),
  1199 => (x"88",x"c1",x"48",x"66"),
  1200 => (x"c5",x"58",x"a6",x"d0"),
  1201 => (x"dc",x"ff",x"87",x"d6"),
  1202 => (x"49",x"70",x"87",x"ce"),
  1203 => (x"59",x"a6",x"ec",x"c0"),
  1204 => (x"87",x"c4",x"dc",x"ff"),
  1205 => (x"e0",x"c0",x"49",x"70"),
  1206 => (x"66",x"dc",x"59",x"a6"),
  1207 => (x"a8",x"ec",x"c0",x"48"),
  1208 => (x"87",x"ca",x"c0",x"05"),
  1209 => (x"c0",x"48",x"a6",x"dc"),
  1210 => (x"c0",x"78",x"66",x"e8"),
  1211 => (x"d8",x"ff",x"87",x"c4"),
  1212 => (x"66",x"c8",x"87",x"f3"),
  1213 => (x"c1",x"91",x"cb",x"49"),
  1214 => (x"71",x"48",x"66",x"c0"),
  1215 => (x"4a",x"7e",x"70",x"80"),
  1216 => (x"49",x"6e",x"82",x"c8"),
  1217 => (x"e8",x"c0",x"81",x"ca"),
  1218 => (x"66",x"dc",x"51",x"66"),
  1219 => (x"c0",x"81",x"c1",x"49"),
  1220 => (x"c1",x"89",x"66",x"e8"),
  1221 => (x"70",x"30",x"71",x"48"),
  1222 => (x"71",x"89",x"c1",x"49"),
  1223 => (x"d1",x"c2",x"7a",x"97"),
  1224 => (x"c0",x"49",x"bf",x"fe"),
  1225 => (x"97",x"29",x"66",x"e8"),
  1226 => (x"71",x"48",x"4a",x"6a"),
  1227 => (x"a6",x"f0",x"c0",x"98"),
  1228 => (x"c4",x"49",x"6e",x"58"),
  1229 => (x"c0",x"4d",x"69",x"81"),
  1230 => (x"c4",x"48",x"66",x"e0"),
  1231 => (x"c0",x"02",x"a8",x"66"),
  1232 => (x"a6",x"c4",x"87",x"c8"),
  1233 => (x"c0",x"78",x"c0",x"48"),
  1234 => (x"a6",x"c4",x"87",x"c5"),
  1235 => (x"c4",x"78",x"c1",x"48"),
  1236 => (x"e0",x"c0",x"1e",x"66"),
  1237 => (x"ff",x"49",x"75",x"1e"),
  1238 => (x"c8",x"87",x"ce",x"d8"),
  1239 => (x"c0",x"4c",x"70",x"86"),
  1240 => (x"c1",x"06",x"ac",x"b7"),
  1241 => (x"85",x"74",x"87",x"d4"),
  1242 => (x"74",x"49",x"e0",x"c0"),
  1243 => (x"c1",x"4b",x"75",x"89"),
  1244 => (x"71",x"4a",x"f7",x"d1"),
  1245 => (x"87",x"ef",x"f4",x"fe"),
  1246 => (x"e4",x"c0",x"85",x"c2"),
  1247 => (x"80",x"c1",x"48",x"66"),
  1248 => (x"58",x"a6",x"e8",x"c0"),
  1249 => (x"49",x"66",x"ec",x"c0"),
  1250 => (x"a9",x"70",x"81",x"c1"),
  1251 => (x"87",x"c8",x"c0",x"02"),
  1252 => (x"c0",x"48",x"a6",x"c4"),
  1253 => (x"87",x"c5",x"c0",x"78"),
  1254 => (x"c1",x"48",x"a6",x"c4"),
  1255 => (x"1e",x"66",x"c4",x"78"),
  1256 => (x"c0",x"49",x"a4",x"c2"),
  1257 => (x"88",x"71",x"48",x"e0"),
  1258 => (x"75",x"1e",x"49",x"70"),
  1259 => (x"f8",x"d6",x"ff",x"49"),
  1260 => (x"c0",x"86",x"c8",x"87"),
  1261 => (x"ff",x"01",x"a8",x"b7"),
  1262 => (x"e4",x"c0",x"87",x"c0"),
  1263 => (x"d1",x"c0",x"02",x"66"),
  1264 => (x"c9",x"49",x"6e",x"87"),
  1265 => (x"66",x"e4",x"c0",x"81"),
  1266 => (x"c0",x"48",x"6e",x"51"),
  1267 => (x"c0",x"78",x"f6",x"fb"),
  1268 => (x"49",x"6e",x"87",x"cc"),
  1269 => (x"51",x"c2",x"81",x"c9"),
  1270 => (x"fd",x"c0",x"48",x"6e"),
  1271 => (x"66",x"c8",x"78",x"e5"),
  1272 => (x"a8",x"66",x"cc",x"48"),
  1273 => (x"87",x"cb",x"c0",x"04"),
  1274 => (x"c1",x"48",x"66",x"c8"),
  1275 => (x"58",x"a6",x"cc",x"80"),
  1276 => (x"cc",x"87",x"e9",x"c0"),
  1277 => (x"88",x"c1",x"48",x"66"),
  1278 => (x"c0",x"58",x"a6",x"d0"),
  1279 => (x"d5",x"ff",x"87",x"de"),
  1280 => (x"4c",x"70",x"87",x"d3"),
  1281 => (x"c1",x"87",x"d5",x"c0"),
  1282 => (x"c0",x"05",x"ac",x"c6"),
  1283 => (x"66",x"d0",x"87",x"c8"),
  1284 => (x"d4",x"80",x"c1",x"48"),
  1285 => (x"d4",x"ff",x"58",x"a6"),
  1286 => (x"4c",x"70",x"87",x"fb"),
  1287 => (x"c1",x"48",x"66",x"d4"),
  1288 => (x"58",x"a6",x"d8",x"80"),
  1289 => (x"c0",x"02",x"9c",x"74"),
  1290 => (x"66",x"c8",x"87",x"cb"),
  1291 => (x"66",x"c8",x"c1",x"48"),
  1292 => (x"e8",x"f2",x"04",x"a8"),
  1293 => (x"d3",x"d4",x"ff",x"87"),
  1294 => (x"48",x"66",x"c8",x"87"),
  1295 => (x"c0",x"03",x"a8",x"c7"),
  1296 => (x"ce",x"c2",x"87",x"e5"),
  1297 => (x"78",x"c0",x"48",x"d2"),
  1298 => (x"cb",x"49",x"66",x"c8"),
  1299 => (x"66",x"c0",x"c1",x"91"),
  1300 => (x"4a",x"a1",x"c4",x"81"),
  1301 => (x"52",x"c0",x"4a",x"6a"),
  1302 => (x"48",x"66",x"c8",x"79"),
  1303 => (x"a6",x"cc",x"80",x"c1"),
  1304 => (x"04",x"a8",x"c7",x"58"),
  1305 => (x"ff",x"87",x"db",x"ff"),
  1306 => (x"de",x"ff",x"8e",x"d0"),
  1307 => (x"6f",x"4c",x"87",x"e5"),
  1308 => (x"2a",x"20",x"64",x"61"),
  1309 => (x"3a",x"00",x"20",x"2e"),
  1310 => (x"73",x"1e",x"00",x"20"),
  1311 => (x"9b",x"4b",x"71",x"1e"),
  1312 => (x"c2",x"87",x"c6",x"02"),
  1313 => (x"c0",x"48",x"ce",x"ce"),
  1314 => (x"c2",x"1e",x"c7",x"78"),
  1315 => (x"49",x"bf",x"ce",x"ce"),
  1316 => (x"cb",x"d3",x"c1",x"1e"),
  1317 => (x"f6",x"cd",x"c2",x"1e"),
  1318 => (x"e8",x"ed",x"49",x"bf"),
  1319 => (x"c2",x"86",x"cc",x"87"),
  1320 => (x"49",x"bf",x"f6",x"cd"),
  1321 => (x"73",x"87",x"e7",x"e8"),
  1322 => (x"87",x"c7",x"02",x"9b"),
  1323 => (x"49",x"cb",x"d3",x"c1"),
  1324 => (x"ff",x"87",x"f3",x"df"),
  1325 => (x"00",x"87",x"e0",x"dd"),
  1326 => (x"00",x"00",x"01",x"00"),
  1327 => (x"45",x"20",x"80",x"00"),
  1328 => (x"00",x"74",x"69",x"78"),
  1329 => (x"61",x"42",x"20",x"80"),
  1330 => (x"69",x"00",x"6b",x"63"),
  1331 => (x"a2",x"00",x"00",x"0c"),
  1332 => (x"00",x"00",x"00",x"23"),
  1333 => (x"0c",x"69",x"00",x"00"),
  1334 => (x"23",x"c0",x"00",x"00"),
  1335 => (x"00",x"00",x"00",x"00"),
  1336 => (x"00",x"0c",x"69",x"00"),
  1337 => (x"00",x"23",x"de",x"00"),
  1338 => (x"00",x"00",x"00",x"00"),
  1339 => (x"00",x"00",x"0c",x"69"),
  1340 => (x"00",x"00",x"23",x"fc"),
  1341 => (x"69",x"00",x"00",x"00"),
  1342 => (x"1a",x"00",x"00",x"0c"),
  1343 => (x"00",x"00",x"00",x"24"),
  1344 => (x"0c",x"69",x"00",x"00"),
  1345 => (x"24",x"38",x"00",x"00"),
  1346 => (x"00",x"00",x"00",x"00"),
  1347 => (x"00",x"0c",x"69",x"00"),
  1348 => (x"00",x"24",x"56",x"00"),
  1349 => (x"00",x"00",x"00",x"00"),
  1350 => (x"00",x"00",x"0e",x"a6"),
  1351 => (x"00",x"00",x"00",x"00"),
  1352 => (x"76",x"00",x"00",x"00"),
  1353 => (x"00",x"00",x"00",x"0f"),
  1354 => (x"00",x"00",x"00",x"00"),
  1355 => (x"fe",x"1e",x"00",x"00"),
  1356 => (x"78",x"c0",x"48",x"f0"),
  1357 => (x"09",x"79",x"09",x"cd"),
  1358 => (x"1e",x"1e",x"4f",x"26"),
  1359 => (x"7e",x"bf",x"f0",x"fe"),
  1360 => (x"4f",x"26",x"26",x"48"),
  1361 => (x"48",x"f0",x"fe",x"1e"),
  1362 => (x"4f",x"26",x"78",x"c1"),
  1363 => (x"48",x"f0",x"fe",x"1e"),
  1364 => (x"4f",x"26",x"78",x"c0"),
  1365 => (x"c0",x"4a",x"71",x"1e"),
  1366 => (x"4f",x"26",x"52",x"52"),
  1367 => (x"5c",x"5b",x"5e",x"0e"),
  1368 => (x"86",x"f4",x"0e",x"5d"),
  1369 => (x"6d",x"97",x"4d",x"71"),
  1370 => (x"4c",x"a5",x"c1",x"7e"),
  1371 => (x"c8",x"48",x"6c",x"97"),
  1372 => (x"48",x"6e",x"58",x"a6"),
  1373 => (x"05",x"a8",x"66",x"c4"),
  1374 => (x"48",x"ff",x"87",x"c5"),
  1375 => (x"ff",x"87",x"e6",x"c0"),
  1376 => (x"a5",x"c2",x"87",x"ca"),
  1377 => (x"4b",x"6c",x"97",x"49"),
  1378 => (x"97",x"4b",x"a3",x"71"),
  1379 => (x"6c",x"97",x"4b",x"6b"),
  1380 => (x"c1",x"48",x"6e",x"7e"),
  1381 => (x"58",x"a6",x"c8",x"80"),
  1382 => (x"a6",x"cc",x"98",x"c7"),
  1383 => (x"7c",x"97",x"70",x"58"),
  1384 => (x"73",x"87",x"e1",x"fe"),
  1385 => (x"26",x"8e",x"f4",x"48"),
  1386 => (x"26",x"4c",x"26",x"4d"),
  1387 => (x"0e",x"4f",x"26",x"4b"),
  1388 => (x"0e",x"5c",x"5b",x"5e"),
  1389 => (x"4c",x"71",x"86",x"f4"),
  1390 => (x"c3",x"4a",x"66",x"d8"),
  1391 => (x"a4",x"c2",x"9a",x"ff"),
  1392 => (x"49",x"6c",x"97",x"4b"),
  1393 => (x"72",x"49",x"a1",x"73"),
  1394 => (x"7e",x"6c",x"97",x"51"),
  1395 => (x"80",x"c1",x"48",x"6e"),
  1396 => (x"c7",x"58",x"a6",x"c8"),
  1397 => (x"58",x"a6",x"cc",x"98"),
  1398 => (x"8e",x"f4",x"54",x"70"),
  1399 => (x"1e",x"87",x"ca",x"ff"),
  1400 => (x"87",x"e8",x"fd",x"1e"),
  1401 => (x"49",x"4a",x"bf",x"e0"),
  1402 => (x"99",x"c0",x"e0",x"c0"),
  1403 => (x"72",x"87",x"cb",x"02"),
  1404 => (x"f4",x"d1",x"c2",x"1e"),
  1405 => (x"87",x"f7",x"fe",x"49"),
  1406 => (x"fd",x"fc",x"86",x"c4"),
  1407 => (x"fd",x"7e",x"70",x"87"),
  1408 => (x"26",x"26",x"87",x"c2"),
  1409 => (x"d1",x"c2",x"1e",x"4f"),
  1410 => (x"c7",x"fd",x"49",x"f4"),
  1411 => (x"df",x"d7",x"c1",x"87"),
  1412 => (x"87",x"da",x"fc",x"49"),
  1413 => (x"26",x"87",x"fe",x"c2"),
  1414 => (x"1e",x"73",x"1e",x"4f"),
  1415 => (x"49",x"f4",x"d1",x"c2"),
  1416 => (x"70",x"87",x"f9",x"fc"),
  1417 => (x"aa",x"b7",x"c0",x"4a"),
  1418 => (x"87",x"cc",x"c2",x"04"),
  1419 => (x"05",x"aa",x"f0",x"c3"),
  1420 => (x"db",x"c1",x"87",x"c9"),
  1421 => (x"78",x"c1",x"48",x"c4"),
  1422 => (x"c3",x"87",x"ed",x"c1"),
  1423 => (x"c9",x"05",x"aa",x"e0"),
  1424 => (x"c8",x"db",x"c1",x"87"),
  1425 => (x"c1",x"78",x"c1",x"48"),
  1426 => (x"db",x"c1",x"87",x"de"),
  1427 => (x"c6",x"02",x"bf",x"c8"),
  1428 => (x"a2",x"c0",x"c2",x"87"),
  1429 => (x"72",x"87",x"c2",x"4b"),
  1430 => (x"c4",x"db",x"c1",x"4b"),
  1431 => (x"e0",x"c0",x"02",x"bf"),
  1432 => (x"c4",x"49",x"73",x"87"),
  1433 => (x"c1",x"91",x"29",x"b7"),
  1434 => (x"73",x"81",x"e4",x"dc"),
  1435 => (x"c2",x"9a",x"cf",x"4a"),
  1436 => (x"72",x"48",x"c1",x"92"),
  1437 => (x"ff",x"4a",x"70",x"30"),
  1438 => (x"69",x"48",x"72",x"ba"),
  1439 => (x"db",x"79",x"70",x"98"),
  1440 => (x"c4",x"49",x"73",x"87"),
  1441 => (x"c1",x"91",x"29",x"b7"),
  1442 => (x"73",x"81",x"e4",x"dc"),
  1443 => (x"c2",x"9a",x"cf",x"4a"),
  1444 => (x"72",x"48",x"c3",x"92"),
  1445 => (x"48",x"4a",x"70",x"30"),
  1446 => (x"79",x"70",x"b0",x"69"),
  1447 => (x"48",x"c8",x"db",x"c1"),
  1448 => (x"db",x"c1",x"78",x"c0"),
  1449 => (x"78",x"c0",x"48",x"c4"),
  1450 => (x"49",x"f4",x"d1",x"c2"),
  1451 => (x"70",x"87",x"ed",x"fa"),
  1452 => (x"aa",x"b7",x"c0",x"4a"),
  1453 => (x"87",x"f4",x"fd",x"03"),
  1454 => (x"87",x"c4",x"48",x"c0"),
  1455 => (x"4c",x"26",x"4d",x"26"),
  1456 => (x"4f",x"26",x"4b",x"26"),
  1457 => (x"00",x"00",x"00",x"00"),
  1458 => (x"00",x"00",x"00",x"00"),
  1459 => (x"49",x"4a",x"71",x"1e"),
  1460 => (x"26",x"87",x"c6",x"fd"),
  1461 => (x"4a",x"c0",x"1e",x"4f"),
  1462 => (x"91",x"c4",x"49",x"72"),
  1463 => (x"81",x"e4",x"dc",x"c1"),
  1464 => (x"82",x"c1",x"79",x"c0"),
  1465 => (x"04",x"aa",x"b7",x"d0"),
  1466 => (x"4f",x"26",x"87",x"ee"),
  1467 => (x"5c",x"5b",x"5e",x"0e"),
  1468 => (x"4d",x"71",x"0e",x"5d"),
  1469 => (x"75",x"87",x"d5",x"f9"),
  1470 => (x"2a",x"b7",x"c4",x"4a"),
  1471 => (x"e4",x"dc",x"c1",x"92"),
  1472 => (x"cf",x"4c",x"75",x"82"),
  1473 => (x"6a",x"94",x"c2",x"9c"),
  1474 => (x"2b",x"74",x"4b",x"49"),
  1475 => (x"48",x"c2",x"9b",x"c3"),
  1476 => (x"4c",x"70",x"30",x"74"),
  1477 => (x"48",x"74",x"bc",x"ff"),
  1478 => (x"7a",x"70",x"98",x"71"),
  1479 => (x"73",x"87",x"e5",x"f8"),
  1480 => (x"87",x"d8",x"fe",x"48"),
  1481 => (x"00",x"00",x"00",x"00"),
  1482 => (x"00",x"00",x"00",x"00"),
  1483 => (x"00",x"00",x"00",x"00"),
  1484 => (x"00",x"00",x"00",x"00"),
  1485 => (x"00",x"00",x"00",x"00"),
  1486 => (x"00",x"00",x"00",x"00"),
  1487 => (x"00",x"00",x"00",x"00"),
  1488 => (x"00",x"00",x"00",x"00"),
  1489 => (x"00",x"00",x"00",x"00"),
  1490 => (x"00",x"00",x"00",x"00"),
  1491 => (x"00",x"00",x"00",x"00"),
  1492 => (x"00",x"00",x"00",x"00"),
  1493 => (x"00",x"00",x"00",x"00"),
  1494 => (x"00",x"00",x"00",x"00"),
  1495 => (x"00",x"00",x"00",x"00"),
  1496 => (x"00",x"00",x"00",x"00"),
  1497 => (x"48",x"d0",x"ff",x"1e"),
  1498 => (x"71",x"78",x"e1",x"c8"),
  1499 => (x"08",x"d4",x"ff",x"48"),
  1500 => (x"48",x"66",x"c4",x"78"),
  1501 => (x"78",x"08",x"d4",x"ff"),
  1502 => (x"71",x"1e",x"4f",x"26"),
  1503 => (x"49",x"66",x"c4",x"4a"),
  1504 => (x"ff",x"49",x"72",x"1e"),
  1505 => (x"d0",x"ff",x"87",x"de"),
  1506 => (x"78",x"e0",x"c0",x"48"),
  1507 => (x"1e",x"4f",x"26",x"26"),
  1508 => (x"4b",x"71",x"1e",x"73"),
  1509 => (x"1e",x"49",x"66",x"c8"),
  1510 => (x"e0",x"c1",x"4a",x"73"),
  1511 => (x"d9",x"ff",x"49",x"a2"),
  1512 => (x"87",x"c4",x"26",x"87"),
  1513 => (x"4c",x"26",x"4d",x"26"),
  1514 => (x"4f",x"26",x"4b",x"26"),
  1515 => (x"71",x"1e",x"73",x"1e"),
  1516 => (x"b7",x"c2",x"4b",x"4a"),
  1517 => (x"87",x"c8",x"03",x"ab"),
  1518 => (x"c3",x"4a",x"49",x"a3"),
  1519 => (x"87",x"c7",x"9a",x"ff"),
  1520 => (x"4a",x"49",x"a3",x"ce"),
  1521 => (x"c8",x"9a",x"ff",x"c3"),
  1522 => (x"72",x"1e",x"49",x"66"),
  1523 => (x"87",x"ea",x"fe",x"49"),
  1524 => (x"87",x"d4",x"ff",x"26"),
  1525 => (x"4a",x"d4",x"ff",x"1e"),
  1526 => (x"ff",x"7a",x"ff",x"c3"),
  1527 => (x"e1",x"c0",x"48",x"d0"),
  1528 => (x"c2",x"7a",x"de",x"78"),
  1529 => (x"7a",x"bf",x"fe",x"d1"),
  1530 => (x"28",x"c8",x"48",x"49"),
  1531 => (x"48",x"71",x"7a",x"70"),
  1532 => (x"7a",x"70",x"28",x"d0"),
  1533 => (x"28",x"d8",x"48",x"71"),
  1534 => (x"d0",x"ff",x"7a",x"70"),
  1535 => (x"78",x"e0",x"c0",x"48"),
  1536 => (x"ff",x"1e",x"4f",x"26"),
  1537 => (x"c9",x"c8",x"48",x"d0"),
  1538 => (x"ff",x"48",x"71",x"78"),
  1539 => (x"26",x"78",x"08",x"d4"),
  1540 => (x"4a",x"71",x"1e",x"4f"),
  1541 => (x"ff",x"87",x"eb",x"49"),
  1542 => (x"78",x"c8",x"48",x"d0"),
  1543 => (x"73",x"1e",x"4f",x"26"),
  1544 => (x"c2",x"4b",x"71",x"1e"),
  1545 => (x"02",x"bf",x"ce",x"d2"),
  1546 => (x"eb",x"c2",x"87",x"c3"),
  1547 => (x"48",x"d0",x"ff",x"87"),
  1548 => (x"73",x"78",x"c9",x"c8"),
  1549 => (x"b1",x"e0",x"c0",x"49"),
  1550 => (x"71",x"48",x"d4",x"ff"),
  1551 => (x"c2",x"d2",x"c2",x"78"),
  1552 => (x"c8",x"78",x"c0",x"48"),
  1553 => (x"87",x"c5",x"02",x"66"),
  1554 => (x"c2",x"49",x"ff",x"c3"),
  1555 => (x"c2",x"49",x"c0",x"87"),
  1556 => (x"cc",x"59",x"ca",x"d2"),
  1557 => (x"87",x"c6",x"02",x"66"),
  1558 => (x"4a",x"d5",x"d5",x"c5"),
  1559 => (x"ff",x"cf",x"87",x"c4"),
  1560 => (x"d2",x"c2",x"4a",x"ff"),
  1561 => (x"d2",x"c2",x"5a",x"ce"),
  1562 => (x"78",x"c1",x"48",x"ce"),
  1563 => (x"4d",x"26",x"87",x"c4"),
  1564 => (x"4b",x"26",x"4c",x"26"),
  1565 => (x"5e",x"0e",x"4f",x"26"),
  1566 => (x"0e",x"5d",x"5c",x"5b"),
  1567 => (x"d2",x"c2",x"4a",x"71"),
  1568 => (x"72",x"4c",x"bf",x"ca"),
  1569 => (x"87",x"cb",x"02",x"9a"),
  1570 => (x"c1",x"91",x"c8",x"49"),
  1571 => (x"71",x"4b",x"d4",x"e0"),
  1572 => (x"c1",x"87",x"c4",x"83"),
  1573 => (x"c0",x"4b",x"d4",x"e4"),
  1574 => (x"74",x"49",x"13",x"4d"),
  1575 => (x"c6",x"d2",x"c2",x"99"),
  1576 => (x"d4",x"ff",x"b9",x"bf"),
  1577 => (x"c1",x"78",x"71",x"48"),
  1578 => (x"c8",x"85",x"2c",x"b7"),
  1579 => (x"e8",x"04",x"ad",x"b7"),
  1580 => (x"c2",x"d2",x"c2",x"87"),
  1581 => (x"80",x"c8",x"48",x"bf"),
  1582 => (x"58",x"c6",x"d2",x"c2"),
  1583 => (x"1e",x"87",x"ef",x"fe"),
  1584 => (x"4b",x"71",x"1e",x"73"),
  1585 => (x"02",x"9a",x"4a",x"13"),
  1586 => (x"49",x"72",x"87",x"cb"),
  1587 => (x"13",x"87",x"e7",x"fe"),
  1588 => (x"f5",x"05",x"9a",x"4a"),
  1589 => (x"87",x"da",x"fe",x"87"),
  1590 => (x"c2",x"d2",x"c2",x"1e"),
  1591 => (x"d2",x"c2",x"49",x"bf"),
  1592 => (x"a1",x"c1",x"48",x"c2"),
  1593 => (x"b7",x"c0",x"c4",x"78"),
  1594 => (x"87",x"db",x"03",x"a9"),
  1595 => (x"c2",x"48",x"d4",x"ff"),
  1596 => (x"78",x"bf",x"c6",x"d2"),
  1597 => (x"bf",x"c2",x"d2",x"c2"),
  1598 => (x"c2",x"d2",x"c2",x"49"),
  1599 => (x"78",x"a1",x"c1",x"48"),
  1600 => (x"a9",x"b7",x"c0",x"c4"),
  1601 => (x"ff",x"87",x"e5",x"04"),
  1602 => (x"78",x"c8",x"48",x"d0"),
  1603 => (x"48",x"ce",x"d2",x"c2"),
  1604 => (x"4f",x"26",x"78",x"c0"),
  1605 => (x"00",x"00",x"00",x"00"),
  1606 => (x"00",x"00",x"00",x"00"),
  1607 => (x"5f",x"00",x"00",x"00"),
  1608 => (x"00",x"00",x"00",x"5f"),
  1609 => (x"00",x"03",x"03",x"00"),
  1610 => (x"00",x"00",x"03",x"03"),
  1611 => (x"14",x"7f",x"7f",x"14"),
  1612 => (x"00",x"14",x"7f",x"7f"),
  1613 => (x"6b",x"2e",x"24",x"00"),
  1614 => (x"00",x"12",x"3a",x"6b"),
  1615 => (x"18",x"36",x"6a",x"4c"),
  1616 => (x"00",x"32",x"56",x"6c"),
  1617 => (x"59",x"4f",x"7e",x"30"),
  1618 => (x"40",x"68",x"3a",x"77"),
  1619 => (x"07",x"04",x"00",x"00"),
  1620 => (x"00",x"00",x"00",x"03"),
  1621 => (x"3e",x"1c",x"00",x"00"),
  1622 => (x"00",x"00",x"41",x"63"),
  1623 => (x"63",x"41",x"00",x"00"),
  1624 => (x"00",x"00",x"1c",x"3e"),
  1625 => (x"1c",x"3e",x"2a",x"08"),
  1626 => (x"08",x"2a",x"3e",x"1c"),
  1627 => (x"3e",x"08",x"08",x"00"),
  1628 => (x"00",x"08",x"08",x"3e"),
  1629 => (x"e0",x"80",x"00",x"00"),
  1630 => (x"00",x"00",x"00",x"60"),
  1631 => (x"08",x"08",x"08",x"00"),
  1632 => (x"00",x"08",x"08",x"08"),
  1633 => (x"60",x"00",x"00",x"00"),
  1634 => (x"00",x"00",x"00",x"60"),
  1635 => (x"18",x"30",x"60",x"40"),
  1636 => (x"01",x"03",x"06",x"0c"),
  1637 => (x"59",x"7f",x"3e",x"00"),
  1638 => (x"00",x"3e",x"7f",x"4d"),
  1639 => (x"7f",x"06",x"04",x"00"),
  1640 => (x"00",x"00",x"00",x"7f"),
  1641 => (x"71",x"63",x"42",x"00"),
  1642 => (x"00",x"46",x"4f",x"59"),
  1643 => (x"49",x"63",x"22",x"00"),
  1644 => (x"00",x"36",x"7f",x"49"),
  1645 => (x"13",x"16",x"1c",x"18"),
  1646 => (x"00",x"10",x"7f",x"7f"),
  1647 => (x"45",x"67",x"27",x"00"),
  1648 => (x"00",x"39",x"7d",x"45"),
  1649 => (x"4b",x"7e",x"3c",x"00"),
  1650 => (x"00",x"30",x"79",x"49"),
  1651 => (x"71",x"01",x"01",x"00"),
  1652 => (x"00",x"07",x"0f",x"79"),
  1653 => (x"49",x"7f",x"36",x"00"),
  1654 => (x"00",x"36",x"7f",x"49"),
  1655 => (x"49",x"4f",x"06",x"00"),
  1656 => (x"00",x"1e",x"3f",x"69"),
  1657 => (x"66",x"00",x"00",x"00"),
  1658 => (x"00",x"00",x"00",x"66"),
  1659 => (x"e6",x"80",x"00",x"00"),
  1660 => (x"00",x"00",x"00",x"66"),
  1661 => (x"14",x"08",x"08",x"00"),
  1662 => (x"00",x"22",x"22",x"14"),
  1663 => (x"14",x"14",x"14",x"00"),
  1664 => (x"00",x"14",x"14",x"14"),
  1665 => (x"14",x"22",x"22",x"00"),
  1666 => (x"00",x"08",x"08",x"14"),
  1667 => (x"51",x"03",x"02",x"00"),
  1668 => (x"00",x"06",x"0f",x"59"),
  1669 => (x"5d",x"41",x"7f",x"3e"),
  1670 => (x"00",x"1e",x"1f",x"55"),
  1671 => (x"09",x"7f",x"7e",x"00"),
  1672 => (x"00",x"7e",x"7f",x"09"),
  1673 => (x"49",x"7f",x"7f",x"00"),
  1674 => (x"00",x"36",x"7f",x"49"),
  1675 => (x"63",x"3e",x"1c",x"00"),
  1676 => (x"00",x"41",x"41",x"41"),
  1677 => (x"41",x"7f",x"7f",x"00"),
  1678 => (x"00",x"1c",x"3e",x"63"),
  1679 => (x"49",x"7f",x"7f",x"00"),
  1680 => (x"00",x"41",x"41",x"49"),
  1681 => (x"09",x"7f",x"7f",x"00"),
  1682 => (x"00",x"01",x"01",x"09"),
  1683 => (x"41",x"7f",x"3e",x"00"),
  1684 => (x"00",x"7a",x"7b",x"49"),
  1685 => (x"08",x"7f",x"7f",x"00"),
  1686 => (x"00",x"7f",x"7f",x"08"),
  1687 => (x"7f",x"41",x"00",x"00"),
  1688 => (x"00",x"00",x"41",x"7f"),
  1689 => (x"40",x"60",x"20",x"00"),
  1690 => (x"00",x"3f",x"7f",x"40"),
  1691 => (x"1c",x"08",x"7f",x"7f"),
  1692 => (x"00",x"41",x"63",x"36"),
  1693 => (x"40",x"7f",x"7f",x"00"),
  1694 => (x"00",x"40",x"40",x"40"),
  1695 => (x"0c",x"06",x"7f",x"7f"),
  1696 => (x"00",x"7f",x"7f",x"06"),
  1697 => (x"0c",x"06",x"7f",x"7f"),
  1698 => (x"00",x"7f",x"7f",x"18"),
  1699 => (x"41",x"7f",x"3e",x"00"),
  1700 => (x"00",x"3e",x"7f",x"41"),
  1701 => (x"09",x"7f",x"7f",x"00"),
  1702 => (x"00",x"06",x"0f",x"09"),
  1703 => (x"61",x"41",x"7f",x"3e"),
  1704 => (x"00",x"40",x"7e",x"7f"),
  1705 => (x"09",x"7f",x"7f",x"00"),
  1706 => (x"00",x"66",x"7f",x"19"),
  1707 => (x"4d",x"6f",x"26",x"00"),
  1708 => (x"00",x"32",x"7b",x"59"),
  1709 => (x"7f",x"01",x"01",x"00"),
  1710 => (x"00",x"01",x"01",x"7f"),
  1711 => (x"40",x"7f",x"3f",x"00"),
  1712 => (x"00",x"3f",x"7f",x"40"),
  1713 => (x"70",x"3f",x"0f",x"00"),
  1714 => (x"00",x"0f",x"3f",x"70"),
  1715 => (x"18",x"30",x"7f",x"7f"),
  1716 => (x"00",x"7f",x"7f",x"30"),
  1717 => (x"1c",x"36",x"63",x"41"),
  1718 => (x"41",x"63",x"36",x"1c"),
  1719 => (x"7c",x"06",x"03",x"01"),
  1720 => (x"01",x"03",x"06",x"7c"),
  1721 => (x"4d",x"59",x"71",x"61"),
  1722 => (x"00",x"41",x"43",x"47"),
  1723 => (x"7f",x"7f",x"00",x"00"),
  1724 => (x"00",x"00",x"41",x"41"),
  1725 => (x"0c",x"06",x"03",x"01"),
  1726 => (x"40",x"60",x"30",x"18"),
  1727 => (x"41",x"41",x"00",x"00"),
  1728 => (x"00",x"00",x"7f",x"7f"),
  1729 => (x"03",x"06",x"0c",x"08"),
  1730 => (x"00",x"08",x"0c",x"06"),
  1731 => (x"80",x"80",x"80",x"80"),
  1732 => (x"00",x"80",x"80",x"80"),
  1733 => (x"03",x"00",x"00",x"00"),
  1734 => (x"00",x"00",x"04",x"07"),
  1735 => (x"54",x"74",x"20",x"00"),
  1736 => (x"00",x"78",x"7c",x"54"),
  1737 => (x"44",x"7f",x"7f",x"00"),
  1738 => (x"00",x"38",x"7c",x"44"),
  1739 => (x"44",x"7c",x"38",x"00"),
  1740 => (x"00",x"00",x"44",x"44"),
  1741 => (x"44",x"7c",x"38",x"00"),
  1742 => (x"00",x"7f",x"7f",x"44"),
  1743 => (x"54",x"7c",x"38",x"00"),
  1744 => (x"00",x"18",x"5c",x"54"),
  1745 => (x"7f",x"7e",x"04",x"00"),
  1746 => (x"00",x"00",x"05",x"05"),
  1747 => (x"a4",x"bc",x"18",x"00"),
  1748 => (x"00",x"7c",x"fc",x"a4"),
  1749 => (x"04",x"7f",x"7f",x"00"),
  1750 => (x"00",x"78",x"7c",x"04"),
  1751 => (x"3d",x"00",x"00",x"00"),
  1752 => (x"00",x"00",x"40",x"7d"),
  1753 => (x"80",x"80",x"80",x"00"),
  1754 => (x"00",x"00",x"7d",x"fd"),
  1755 => (x"10",x"7f",x"7f",x"00"),
  1756 => (x"00",x"44",x"6c",x"38"),
  1757 => (x"3f",x"00",x"00",x"00"),
  1758 => (x"00",x"00",x"40",x"7f"),
  1759 => (x"18",x"0c",x"7c",x"7c"),
  1760 => (x"00",x"78",x"7c",x"0c"),
  1761 => (x"04",x"7c",x"7c",x"00"),
  1762 => (x"00",x"78",x"7c",x"04"),
  1763 => (x"44",x"7c",x"38",x"00"),
  1764 => (x"00",x"38",x"7c",x"44"),
  1765 => (x"24",x"fc",x"fc",x"00"),
  1766 => (x"00",x"18",x"3c",x"24"),
  1767 => (x"24",x"3c",x"18",x"00"),
  1768 => (x"00",x"fc",x"fc",x"24"),
  1769 => (x"04",x"7c",x"7c",x"00"),
  1770 => (x"00",x"08",x"0c",x"04"),
  1771 => (x"54",x"5c",x"48",x"00"),
  1772 => (x"00",x"20",x"74",x"54"),
  1773 => (x"7f",x"3f",x"04",x"00"),
  1774 => (x"00",x"00",x"44",x"44"),
  1775 => (x"40",x"7c",x"3c",x"00"),
  1776 => (x"00",x"7c",x"7c",x"40"),
  1777 => (x"60",x"3c",x"1c",x"00"),
  1778 => (x"00",x"1c",x"3c",x"60"),
  1779 => (x"30",x"60",x"7c",x"3c"),
  1780 => (x"00",x"3c",x"7c",x"60"),
  1781 => (x"10",x"38",x"6c",x"44"),
  1782 => (x"00",x"44",x"6c",x"38"),
  1783 => (x"e0",x"bc",x"1c",x"00"),
  1784 => (x"00",x"1c",x"3c",x"60"),
  1785 => (x"74",x"64",x"44",x"00"),
  1786 => (x"00",x"44",x"4c",x"5c"),
  1787 => (x"3e",x"08",x"08",x"00"),
  1788 => (x"00",x"41",x"41",x"77"),
  1789 => (x"7f",x"00",x"00",x"00"),
  1790 => (x"00",x"00",x"00",x"7f"),
  1791 => (x"77",x"41",x"41",x"00"),
  1792 => (x"00",x"08",x"08",x"3e"),
  1793 => (x"03",x"01",x"01",x"02"),
  1794 => (x"00",x"01",x"02",x"02"),
  1795 => (x"7f",x"7f",x"7f",x"7f"),
  1796 => (x"00",x"7f",x"7f",x"7f"),
  1797 => (x"1c",x"1c",x"08",x"08"),
  1798 => (x"7f",x"7f",x"3e",x"3e"),
  1799 => (x"3e",x"3e",x"7f",x"7f"),
  1800 => (x"08",x"08",x"1c",x"1c"),
  1801 => (x"7c",x"18",x"10",x"00"),
  1802 => (x"00",x"10",x"18",x"7c"),
  1803 => (x"7c",x"30",x"10",x"00"),
  1804 => (x"00",x"10",x"30",x"7c"),
  1805 => (x"60",x"60",x"30",x"10"),
  1806 => (x"00",x"06",x"1e",x"78"),
  1807 => (x"18",x"3c",x"66",x"42"),
  1808 => (x"00",x"42",x"66",x"3c"),
  1809 => (x"c2",x"6a",x"38",x"78"),
  1810 => (x"00",x"38",x"6c",x"c6"),
  1811 => (x"60",x"00",x"00",x"60"),
  1812 => (x"00",x"60",x"00",x"00"),
  1813 => (x"5c",x"5b",x"5e",x"0e"),
  1814 => (x"71",x"1e",x"0e",x"5d"),
  1815 => (x"df",x"d2",x"c2",x"4c"),
  1816 => (x"4b",x"c0",x"4d",x"bf"),
  1817 => (x"ab",x"74",x"1e",x"c0"),
  1818 => (x"c4",x"87",x"c7",x"02"),
  1819 => (x"78",x"c0",x"48",x"a6"),
  1820 => (x"a6",x"c4",x"87",x"c5"),
  1821 => (x"c4",x"78",x"c1",x"48"),
  1822 => (x"49",x"73",x"1e",x"66"),
  1823 => (x"c8",x"87",x"df",x"ee"),
  1824 => (x"49",x"e0",x"c0",x"86"),
  1825 => (x"c4",x"87",x"ef",x"ef"),
  1826 => (x"49",x"6a",x"4a",x"a5"),
  1827 => (x"f1",x"87",x"f0",x"f0"),
  1828 => (x"85",x"cb",x"87",x"c6"),
  1829 => (x"b7",x"c8",x"83",x"c1"),
  1830 => (x"c7",x"ff",x"04",x"ab"),
  1831 => (x"4d",x"26",x"26",x"87"),
  1832 => (x"4b",x"26",x"4c",x"26"),
  1833 => (x"71",x"1e",x"4f",x"26"),
  1834 => (x"e3",x"d2",x"c2",x"4a"),
  1835 => (x"e3",x"d2",x"c2",x"5a"),
  1836 => (x"49",x"78",x"c7",x"48"),
  1837 => (x"26",x"87",x"dd",x"fe"),
  1838 => (x"1e",x"73",x"1e",x"4f"),
  1839 => (x"b7",x"c0",x"4a",x"71"),
  1840 => (x"87",x"d3",x"03",x"aa"),
  1841 => (x"bf",x"e6",x"ff",x"c1"),
  1842 => (x"c1",x"87",x"c4",x"05"),
  1843 => (x"c0",x"87",x"c2",x"4b"),
  1844 => (x"ea",x"ff",x"c1",x"4b"),
  1845 => (x"c1",x"87",x"c4",x"5b"),
  1846 => (x"c1",x"5a",x"ea",x"ff"),
  1847 => (x"4a",x"bf",x"e6",x"ff"),
  1848 => (x"c0",x"c1",x"9a",x"c1"),
  1849 => (x"e8",x"ec",x"49",x"a2"),
  1850 => (x"c1",x"48",x"fc",x"87"),
  1851 => (x"78",x"bf",x"e6",x"ff"),
  1852 => (x"1e",x"87",x"ef",x"fe"),
  1853 => (x"66",x"c4",x"4a",x"71"),
  1854 => (x"ea",x"49",x"72",x"1e"),
  1855 => (x"26",x"26",x"87",x"ee"),
  1856 => (x"4a",x"71",x"1e",x"4f"),
  1857 => (x"c3",x"48",x"d4",x"ff"),
  1858 => (x"d0",x"ff",x"78",x"ff"),
  1859 => (x"78",x"e1",x"c0",x"48"),
  1860 => (x"c1",x"48",x"d4",x"ff"),
  1861 => (x"c4",x"49",x"72",x"78"),
  1862 => (x"ff",x"78",x"71",x"31"),
  1863 => (x"e0",x"c0",x"48",x"d0"),
  1864 => (x"1e",x"4f",x"26",x"78"),
  1865 => (x"bf",x"e6",x"ff",x"c1"),
  1866 => (x"87",x"e0",x"e6",x"49"),
  1867 => (x"48",x"d7",x"d2",x"c2"),
  1868 => (x"c2",x"78",x"bf",x"e8"),
  1869 => (x"ec",x"48",x"d3",x"d2"),
  1870 => (x"d2",x"c2",x"78",x"bf"),
  1871 => (x"49",x"4a",x"bf",x"d7"),
  1872 => (x"c8",x"99",x"ff",x"c3"),
  1873 => (x"48",x"72",x"2a",x"b7"),
  1874 => (x"d2",x"c2",x"b0",x"71"),
  1875 => (x"4f",x"26",x"58",x"df"),
  1876 => (x"5c",x"5b",x"5e",x"0e"),
  1877 => (x"4b",x"71",x"0e",x"5d"),
  1878 => (x"c2",x"87",x"c8",x"ff"),
  1879 => (x"c0",x"48",x"d2",x"d2"),
  1880 => (x"e6",x"49",x"73",x"50"),
  1881 => (x"49",x"70",x"87",x"c6"),
  1882 => (x"cb",x"9c",x"c2",x"4c"),
  1883 => (x"fd",x"c9",x"49",x"ee"),
  1884 => (x"4d",x"49",x"70",x"87"),
  1885 => (x"97",x"d2",x"d2",x"c2"),
  1886 => (x"e2",x"c1",x"05",x"bf"),
  1887 => (x"49",x"66",x"d0",x"87"),
  1888 => (x"bf",x"db",x"d2",x"c2"),
  1889 => (x"87",x"d6",x"05",x"99"),
  1890 => (x"c2",x"49",x"66",x"d4"),
  1891 => (x"99",x"bf",x"d3",x"d2"),
  1892 => (x"73",x"87",x"cb",x"05"),
  1893 => (x"87",x"d4",x"e5",x"49"),
  1894 => (x"c1",x"02",x"98",x"70"),
  1895 => (x"4c",x"c1",x"87",x"c1"),
  1896 => (x"75",x"87",x"c0",x"fe"),
  1897 => (x"87",x"d2",x"c9",x"49"),
  1898 => (x"c6",x"02",x"98",x"70"),
  1899 => (x"d2",x"d2",x"c2",x"87"),
  1900 => (x"c2",x"50",x"c1",x"48"),
  1901 => (x"bf",x"97",x"d2",x"d2"),
  1902 => (x"87",x"e3",x"c0",x"05"),
  1903 => (x"bf",x"db",x"d2",x"c2"),
  1904 => (x"99",x"66",x"d0",x"49"),
  1905 => (x"87",x"d6",x"ff",x"05"),
  1906 => (x"bf",x"d3",x"d2",x"c2"),
  1907 => (x"99",x"66",x"d4",x"49"),
  1908 => (x"87",x"ca",x"ff",x"05"),
  1909 => (x"d3",x"e4",x"49",x"73"),
  1910 => (x"05",x"98",x"70",x"87"),
  1911 => (x"74",x"87",x"ff",x"fe"),
  1912 => (x"87",x"fa",x"fa",x"48"),
  1913 => (x"5c",x"5b",x"5e",x"0e"),
  1914 => (x"86",x"f8",x"0e",x"5d"),
  1915 => (x"ec",x"4c",x"4d",x"c0"),
  1916 => (x"a6",x"c4",x"7e",x"bf"),
  1917 => (x"df",x"d2",x"c2",x"48"),
  1918 => (x"1e",x"c1",x"78",x"bf"),
  1919 => (x"49",x"c7",x"1e",x"c0"),
  1920 => (x"c8",x"87",x"cd",x"fd"),
  1921 => (x"02",x"98",x"70",x"86"),
  1922 => (x"49",x"ff",x"87",x"cd"),
  1923 => (x"c1",x"87",x"ea",x"fa"),
  1924 => (x"d7",x"e3",x"49",x"da"),
  1925 => (x"c2",x"4d",x"c1",x"87"),
  1926 => (x"bf",x"97",x"d2",x"d2"),
  1927 => (x"c1",x"87",x"cf",x"02"),
  1928 => (x"49",x"bf",x"de",x"ff"),
  1929 => (x"ff",x"c1",x"b9",x"c1"),
  1930 => (x"fb",x"71",x"59",x"e2"),
  1931 => (x"d2",x"c2",x"87",x"d3"),
  1932 => (x"c1",x"4b",x"bf",x"d7"),
  1933 => (x"05",x"bf",x"e6",x"ff"),
  1934 => (x"c3",x"87",x"e9",x"c0"),
  1935 => (x"eb",x"e2",x"49",x"fd"),
  1936 => (x"49",x"fa",x"c3",x"87"),
  1937 => (x"73",x"87",x"e5",x"e2"),
  1938 => (x"99",x"ff",x"c3",x"49"),
  1939 => (x"49",x"c0",x"1e",x"71"),
  1940 => (x"73",x"87",x"e0",x"fa"),
  1941 => (x"29",x"b7",x"c8",x"49"),
  1942 => (x"49",x"c1",x"1e",x"71"),
  1943 => (x"c8",x"87",x"d4",x"fa"),
  1944 => (x"87",x"f5",x"c5",x"86"),
  1945 => (x"bf",x"db",x"d2",x"c2"),
  1946 => (x"dd",x"02",x"9b",x"4b"),
  1947 => (x"e2",x"ff",x"c1",x"87"),
  1948 => (x"c5",x"c6",x"49",x"bf"),
  1949 => (x"05",x"98",x"70",x"87"),
  1950 => (x"4b",x"c0",x"87",x"c4"),
  1951 => (x"e0",x"c2",x"87",x"d2"),
  1952 => (x"87",x"ea",x"c5",x"49"),
  1953 => (x"58",x"e6",x"ff",x"c1"),
  1954 => (x"ff",x"c1",x"87",x"c6"),
  1955 => (x"78",x"c0",x"48",x"e2"),
  1956 => (x"99",x"c2",x"49",x"73"),
  1957 => (x"c3",x"87",x"cd",x"05"),
  1958 => (x"cf",x"e1",x"49",x"eb"),
  1959 => (x"c2",x"49",x"70",x"87"),
  1960 => (x"87",x"c2",x"02",x"99"),
  1961 => (x"49",x"73",x"4c",x"fb"),
  1962 => (x"cd",x"05",x"99",x"c1"),
  1963 => (x"49",x"f4",x"c3",x"87"),
  1964 => (x"70",x"87",x"f9",x"e0"),
  1965 => (x"02",x"99",x"c2",x"49"),
  1966 => (x"4c",x"fa",x"87",x"c2"),
  1967 => (x"99",x"c8",x"49",x"73"),
  1968 => (x"c3",x"87",x"cd",x"05"),
  1969 => (x"e3",x"e0",x"49",x"f5"),
  1970 => (x"c2",x"49",x"70",x"87"),
  1971 => (x"87",x"d5",x"02",x"99"),
  1972 => (x"bf",x"e3",x"d2",x"c2"),
  1973 => (x"48",x"87",x"ca",x"02"),
  1974 => (x"d2",x"c2",x"88",x"c1"),
  1975 => (x"c2",x"c0",x"58",x"e7"),
  1976 => (x"c1",x"4c",x"ff",x"87"),
  1977 => (x"c4",x"49",x"73",x"4d"),
  1978 => (x"87",x"ce",x"05",x"99"),
  1979 => (x"ff",x"49",x"f2",x"c3"),
  1980 => (x"70",x"87",x"f9",x"df"),
  1981 => (x"02",x"99",x"c2",x"49"),
  1982 => (x"d2",x"c2",x"87",x"dc"),
  1983 => (x"48",x"7e",x"bf",x"e3"),
  1984 => (x"03",x"a8",x"b7",x"c7"),
  1985 => (x"6e",x"87",x"cb",x"c0"),
  1986 => (x"c2",x"80",x"c1",x"48"),
  1987 => (x"c0",x"58",x"e7",x"d2"),
  1988 => (x"4c",x"fe",x"87",x"c2"),
  1989 => (x"fd",x"c3",x"4d",x"c1"),
  1990 => (x"cf",x"df",x"ff",x"49"),
  1991 => (x"c2",x"49",x"70",x"87"),
  1992 => (x"87",x"d5",x"02",x"99"),
  1993 => (x"bf",x"e3",x"d2",x"c2"),
  1994 => (x"87",x"c9",x"c0",x"02"),
  1995 => (x"48",x"e3",x"d2",x"c2"),
  1996 => (x"c2",x"c0",x"78",x"c0"),
  1997 => (x"c1",x"4c",x"fd",x"87"),
  1998 => (x"49",x"fa",x"c3",x"4d"),
  1999 => (x"87",x"ec",x"de",x"ff"),
  2000 => (x"99",x"c2",x"49",x"70"),
  2001 => (x"87",x"d9",x"c0",x"02"),
  2002 => (x"bf",x"e3",x"d2",x"c2"),
  2003 => (x"a8",x"b7",x"c7",x"48"),
  2004 => (x"87",x"c9",x"c0",x"03"),
  2005 => (x"48",x"e3",x"d2",x"c2"),
  2006 => (x"c2",x"c0",x"78",x"c7"),
  2007 => (x"c1",x"4c",x"fc",x"87"),
  2008 => (x"ac",x"b7",x"c0",x"4d"),
  2009 => (x"87",x"d3",x"c0",x"03"),
  2010 => (x"c1",x"48",x"66",x"c4"),
  2011 => (x"7e",x"70",x"80",x"d8"),
  2012 => (x"c0",x"02",x"bf",x"6e"),
  2013 => (x"74",x"4b",x"87",x"c5"),
  2014 => (x"c0",x"0f",x"73",x"49"),
  2015 => (x"1e",x"f0",x"c3",x"1e"),
  2016 => (x"f7",x"49",x"da",x"c1"),
  2017 => (x"86",x"c8",x"87",x"ca"),
  2018 => (x"c0",x"02",x"98",x"70"),
  2019 => (x"d2",x"c2",x"87",x"d8"),
  2020 => (x"6e",x"7e",x"bf",x"e3"),
  2021 => (x"c4",x"91",x"cb",x"49"),
  2022 => (x"82",x"71",x"4a",x"66"),
  2023 => (x"c5",x"c0",x"02",x"6a"),
  2024 => (x"49",x"6e",x"4b",x"87"),
  2025 => (x"9d",x"75",x"0f",x"73"),
  2026 => (x"87",x"c8",x"c0",x"02"),
  2027 => (x"bf",x"e3",x"d2",x"c2"),
  2028 => (x"87",x"e0",x"f2",x"49"),
  2029 => (x"bf",x"ea",x"ff",x"c1"),
  2030 => (x"87",x"dd",x"c0",x"02"),
  2031 => (x"87",x"fa",x"c0",x"49"),
  2032 => (x"c0",x"02",x"98",x"70"),
  2033 => (x"d2",x"c2",x"87",x"d3"),
  2034 => (x"f2",x"49",x"bf",x"e3"),
  2035 => (x"49",x"c0",x"87",x"c6"),
  2036 => (x"c1",x"87",x"e6",x"f3"),
  2037 => (x"c0",x"48",x"ea",x"ff"),
  2038 => (x"f3",x"8e",x"f8",x"78"),
  2039 => (x"00",x"00",x"87",x"c0"),
  2040 => (x"00",x"00",x"00",x"00"),
  2041 => (x"00",x"00",x"00",x"00"),
  2042 => (x"00",x"00",x"00",x"00"),
  2043 => (x"71",x"1e",x"00",x"00"),
  2044 => (x"bf",x"c8",x"ff",x"4a"),
  2045 => (x"48",x"a1",x"72",x"49"),
  2046 => (x"ff",x"1e",x"4f",x"26"),
  2047 => (x"fe",x"89",x"bf",x"c8"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

