library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"e8d2c287",
    12 => x"86c0c84e",
    13 => x"49e8d2c2",
    14 => x"48f4c0c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087c8ff",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d60299",
    50 => x"c348d4ff",
    51 => x"526878ff",
    52 => x"484966c4",
    53 => x"a6c888c1",
    54 => x"05997158",
    55 => x"4f2687ea",
    56 => x"ff1e731e",
    57 => x"ffc34bd4",
    58 => x"c34a6b7b",
    59 => x"496b7bff",
    60 => x"b17232c8",
    61 => x"6b7bffc3",
    62 => x"7131c84a",
    63 => x"7bffc3b2",
    64 => x"32c8496b",
    65 => x"4871b172",
    66 => x"4d2687c4",
    67 => x"4b264c26",
    68 => x"5e0e4f26",
    69 => x"0e5d5c5b",
    70 => x"d4ff4a71",
    71 => x"c349724c",
    72 => x"7c7199ff",
    73 => x"bff4c0c2",
    74 => x"d087c805",
    75 => x"30c94866",
    76 => x"d058a6d4",
    77 => x"29d84966",
    78 => x"7199ffc3",
    79 => x"4966d07c",
    80 => x"ffc329d0",
    81 => x"d07c7199",
    82 => x"29c84966",
    83 => x"7199ffc3",
    84 => x"4966d07c",
    85 => x"7199ffc3",
    86 => x"d049727c",
    87 => x"99ffc329",
    88 => x"4b6c7c71",
    89 => x"4dfff0c9",
    90 => x"05abffc3",
    91 => x"ffc387d0",
    92 => x"c14b6c7c",
    93 => x"87c6028d",
    94 => x"02abffc3",
    95 => x"487387f0",
    96 => x"0e87c7fe",
    97 => x"5d5c5b5e",
    98 => x"c04b710e",
    99 => x"cdeec54c",
   100 => x"d4ff4adf",
   101 => x"78ffc348",
   102 => x"fec34968",
   103 => x"fdc005a9",
   104 => x"734d7087",
   105 => x"87cc029b",
   106 => x"731e66d0",
   107 => x"87c7fc49",
   108 => x"87d686c4",
   109 => x"c448d0ff",
   110 => x"ffc378d1",
   111 => x"4866d07d",
   112 => x"a6d488c1",
   113 => x"05987058",
   114 => x"d4ff87f0",
   115 => x"78ffc348",
   116 => x"059b7378",
   117 => x"d0ff87c5",
   118 => x"c178d048",
   119 => x"8ac14c4a",
   120 => x"87eefe05",
   121 => x"e1fc4874",
   122 => x"1e731e87",
   123 => x"4bc04a71",
   124 => x"c348d4ff",
   125 => x"d0ff78ff",
   126 => x"78c3c448",
   127 => x"c348d4ff",
   128 => x"1e7278ff",
   129 => x"c1f0ffc0",
   130 => x"c5fc49d1",
   131 => x"7086c487",
   132 => x"87d20598",
   133 => x"cc1ec0c8",
   134 => x"e6fd4966",
   135 => x"7086c487",
   136 => x"48d0ff4b",
   137 => x"487378c2",
   138 => x"0e87e3fb",
   139 => x"5d5c5b5e",
   140 => x"c286f80e",
   141 => x"c048ccc9",
   142 => x"c4c1c278",
   143 => x"fe49c01e",
   144 => x"86c487e7",
   145 => x"c5059870",
   146 => x"c948c087",
   147 => x"4dc087cc",
   148 => x"e4c07ec1",
   149 => x"c249bfcf",
   150 => x"714afac1",
   151 => x"c8f84bc8",
   152 => x"05987087",
   153 => x"7ec087c2",
   154 => x"bfcbe4c0",
   155 => x"d6c2c249",
   156 => x"4bc8714a",
   157 => x"7087f2f7",
   158 => x"87c20598",
   159 => x"026e7ec0",
   160 => x"c287fdc0",
   161 => x"4dbfcac8",
   162 => x"9fc2c9c2",
   163 => x"c5487ebf",
   164 => x"05a8ead6",
   165 => x"c8c287c7",
   166 => x"ce4dbfca",
   167 => x"ca486e87",
   168 => x"02a8d5e9",
   169 => x"48c087c5",
   170 => x"c287efc7",
   171 => x"751ec4c1",
   172 => x"87f5fc49",
   173 => x"987086c4",
   174 => x"c087c505",
   175 => x"87dac748",
   176 => x"bfcbe4c0",
   177 => x"d6c2c249",
   178 => x"4bc8714a",
   179 => x"7087daf6",
   180 => x"87c80598",
   181 => x"48ccc9c2",
   182 => x"87d978c1",
   183 => x"bfcfe4c0",
   184 => x"fac1c249",
   185 => x"4bc8714a",
   186 => x"7087fef5",
   187 => x"87c50298",
   188 => x"e5c648c0",
   189 => x"c2c9c287",
   190 => x"c149bf97",
   191 => x"cd05a9d5",
   192 => x"c3c9c287",
   193 => x"c249bf97",
   194 => x"c002a9ea",
   195 => x"48c087c5",
   196 => x"c287c7c6",
   197 => x"bf97c4c1",
   198 => x"e9c3487e",
   199 => x"cec002a8",
   200 => x"c3486e87",
   201 => x"c002a8eb",
   202 => x"48c087c5",
   203 => x"c287ebc5",
   204 => x"bf97cfc1",
   205 => x"c0059949",
   206 => x"c1c287cc",
   207 => x"49bf97d0",
   208 => x"c002a9c2",
   209 => x"48c087c5",
   210 => x"c287cfc5",
   211 => x"bf97d1c1",
   212 => x"c8c9c248",
   213 => x"484c7058",
   214 => x"c9c288c1",
   215 => x"c1c258cc",
   216 => x"49bf97d2",
   217 => x"c1c28175",
   218 => x"4abf97d3",
   219 => x"a17232c8",
   220 => x"d9cdc27e",
   221 => x"c2786e48",
   222 => x"bf97d4c1",
   223 => x"58a6c848",
   224 => x"bfccc9c2",
   225 => x"87d4c202",
   226 => x"bfcbe4c0",
   227 => x"d6c2c249",
   228 => x"4bc8714a",
   229 => x"7087d2f3",
   230 => x"c5c00298",
   231 => x"c348c087",
   232 => x"c9c287f8",
   233 => x"c24cbfc4",
   234 => x"c25cedcd",
   235 => x"bf97e9c1",
   236 => x"c231c849",
   237 => x"bf97e8c1",
   238 => x"c249a14a",
   239 => x"bf97eac1",
   240 => x"7232d04a",
   241 => x"c1c249a1",
   242 => x"4abf97eb",
   243 => x"a17232d8",
   244 => x"9166c449",
   245 => x"bfd9cdc2",
   246 => x"e1cdc281",
   247 => x"f1c1c259",
   248 => x"c84abf97",
   249 => x"f0c1c232",
   250 => x"a24bbf97",
   251 => x"f2c1c24a",
   252 => x"d04bbf97",
   253 => x"4aa27333",
   254 => x"97f3c1c2",
   255 => x"9bcf4bbf",
   256 => x"a27333d8",
   257 => x"e5cdc24a",
   258 => x"e1cdc25a",
   259 => x"8ac24abf",
   260 => x"cdc29274",
   261 => x"a17248e5",
   262 => x"87cac178",
   263 => x"97d6c1c2",
   264 => x"31c849bf",
   265 => x"97d5c1c2",
   266 => x"49a14abf",
   267 => x"59d4c9c2",
   268 => x"bfd0c9c2",
   269 => x"c731c549",
   270 => x"29c981ff",
   271 => x"59edcdc2",
   272 => x"97dbc1c2",
   273 => x"32c84abf",
   274 => x"97dac1c2",
   275 => x"4aa24bbf",
   276 => x"6e9266c4",
   277 => x"e9cdc282",
   278 => x"e1cdc25a",
   279 => x"c278c048",
   280 => x"7248ddcd",
   281 => x"cdc278a1",
   282 => x"cdc248ed",
   283 => x"c278bfe1",
   284 => x"c248f1cd",
   285 => x"78bfe5cd",
   286 => x"bfccc9c2",
   287 => x"87c9c002",
   288 => x"30c44874",
   289 => x"c9c07e70",
   290 => x"e9cdc287",
   291 => x"30c448bf",
   292 => x"c9c27e70",
   293 => x"786e48d0",
   294 => x"8ef848c1",
   295 => x"4c264d26",
   296 => x"4f264b26",
   297 => x"5c5b5e0e",
   298 => x"4a710e5d",
   299 => x"bfccc9c2",
   300 => x"7287cb02",
   301 => x"722bc74b",
   302 => x"9cffc14c",
   303 => x"4b7287c9",
   304 => x"4c722bc8",
   305 => x"c29cffc3",
   306 => x"83bfd9cd",
   307 => x"bfc7e4c0",
   308 => x"87d902ab",
   309 => x"5bcbe4c0",
   310 => x"1ec4c1c2",
   311 => x"c8f44973",
   312 => x"7086c487",
   313 => x"87c50598",
   314 => x"e6c048c0",
   315 => x"ccc9c287",
   316 => x"87d202bf",
   317 => x"91c44974",
   318 => x"81c4c1c2",
   319 => x"ffcf4d69",
   320 => x"9dffffff",
   321 => x"497487cb",
   322 => x"c1c291c2",
   323 => x"699f81c4",
   324 => x"fe48754d",
   325 => x"5e0e87c6",
   326 => x"0e5d5c5b",
   327 => x"4c7186f8",
   328 => x"87c5059c",
   329 => x"c1c348c0",
   330 => x"7ea4c887",
   331 => x"d878c048",
   332 => x"87c70266",
   333 => x"bf9766d8",
   334 => x"c087c505",
   335 => x"87eac248",
   336 => x"49c11ec0",
   337 => x"87e6c749",
   338 => x"4d7086c4",
   339 => x"c2c1029d",
   340 => x"d4c9c287",
   341 => x"4966d84a",
   342 => x"7087f3eb",
   343 => x"f2c00298",
   344 => x"d84a7587",
   345 => x"4bcb4966",
   346 => x"7087d8ec",
   347 => x"e2c00298",
   348 => x"751ec087",
   349 => x"87c7029d",
   350 => x"c048a6c8",
   351 => x"c887c578",
   352 => x"78c148a6",
   353 => x"c64966c8",
   354 => x"86c487e4",
   355 => x"059d4d70",
   356 => x"7587fefe",
   357 => x"cfc1029d",
   358 => x"49a5dc87",
   359 => x"7869486e",
   360 => x"c449a5da",
   361 => x"a4c448a6",
   362 => x"48699f78",
   363 => x"780866c4",
   364 => x"bfccc9c2",
   365 => x"d487d202",
   366 => x"699f49a5",
   367 => x"ffffc049",
   368 => x"d0487199",
   369 => x"c27e7030",
   370 => x"6e7ec087",
   371 => x"66c44849",
   372 => x"66c480bf",
   373 => x"7cc07808",
   374 => x"c449a4cc",
   375 => x"d079bf66",
   376 => x"79c049a4",
   377 => x"87c248c1",
   378 => x"8ef848c0",
   379 => x"0e87edfa",
   380 => x"5d5c5b5e",
   381 => x"9c4c710e",
   382 => x"87cac102",
   383 => x"6949a4c8",
   384 => x"87c2c102",
   385 => x"6c4a66d0",
   386 => x"a6d48249",
   387 => x"4d66d05a",
   388 => x"c8c9c2b9",
   389 => x"baff4abf",
   390 => x"99719972",
   391 => x"87e4c002",
   392 => x"6b4ba4c4",
   393 => x"87fcf949",
   394 => x"c9c27b70",
   395 => x"6c49bfc4",
   396 => x"757c7181",
   397 => x"c8c9c2b9",
   398 => x"baff4abf",
   399 => x"99719972",
   400 => x"87dcff05",
   401 => x"d3f97c75",
   402 => x"1e731e87",
   403 => x"029b4b71",
   404 => x"a3c887c7",
   405 => x"c5056949",
   406 => x"c048c087",
   407 => x"cdc287f7",
   408 => x"c44abfdd",
   409 => x"496949a3",
   410 => x"c9c289c2",
   411 => x"7191bfc4",
   412 => x"c9c24aa2",
   413 => x"6b49bfc8",
   414 => x"4aa27199",
   415 => x"5acbe4c0",
   416 => x"721e66c8",
   417 => x"87e1ed49",
   418 => x"987086c4",
   419 => x"c087c405",
   420 => x"c187c248",
   421 => x"87c8f848",
   422 => x"711e731e",
   423 => x"c0029b4b",
   424 => x"cdc287e4",
   425 => x"4a735bf1",
   426 => x"c9c28ac2",
   427 => x"9249bfc4",
   428 => x"bfddcdc2",
   429 => x"c2807248",
   430 => x"7158f5cd",
   431 => x"c230c448",
   432 => x"c058d4c9",
   433 => x"cdc287ed",
   434 => x"cdc248ed",
   435 => x"c278bfe1",
   436 => x"c248f1cd",
   437 => x"78bfe5cd",
   438 => x"bfccc9c2",
   439 => x"c287c902",
   440 => x"49bfc4c9",
   441 => x"87c731c4",
   442 => x"bfe9cdc2",
   443 => x"c231c449",
   444 => x"f659d4c9",
   445 => x"5e0e87ea",
   446 => x"710e5c5b",
   447 => x"724bc04a",
   448 => x"e1c0029a",
   449 => x"49a2da87",
   450 => x"c24b699f",
   451 => x"02bfccc9",
   452 => x"a2d487cf",
   453 => x"49699f49",
   454 => x"ffffc04c",
   455 => x"c234d09c",
   456 => x"744cc087",
   457 => x"4973b349",
   458 => x"f587edfd",
   459 => x"5e0e87f0",
   460 => x"0e5d5c5b",
   461 => x"4a7186f4",
   462 => x"9a727ec0",
   463 => x"c287d802",
   464 => x"c048c0c1",
   465 => x"f8c0c278",
   466 => x"f1cdc248",
   467 => x"c0c278bf",
   468 => x"cdc248fc",
   469 => x"c278bfed",
   470 => x"c048e1c9",
   471 => x"d0c9c250",
   472 => x"c1c249bf",
   473 => x"714abfc0",
   474 => x"c7c403aa",
   475 => x"cf497287",
   476 => x"e9c00599",
   477 => x"c7e4c087",
   478 => x"f8c0c248",
   479 => x"c1c278bf",
   480 => x"c0c21ec4",
   481 => x"c249bff8",
   482 => x"c148f8c0",
   483 => x"e97178a1",
   484 => x"86c487d7",
   485 => x"48c3e4c0",
   486 => x"78c4c1c2",
   487 => x"e4c087cc",
   488 => x"c048bfc3",
   489 => x"e4c080e0",
   490 => x"c1c258c7",
   491 => x"c148bfc0",
   492 => x"c4c1c280",
   493 => x"09032758",
   494 => x"97bf0000",
   495 => x"029d4dbf",
   496 => x"c387e1c2",
   497 => x"c202ade5",
   498 => x"e4c087da",
   499 => x"cb4bbfc3",
   500 => x"4c1149a3",
   501 => x"c105accf",
   502 => x"497587d2",
   503 => x"89c199df",
   504 => x"c9c291cd",
   505 => x"a3c181d4",
   506 => x"c351124a",
   507 => x"51124aa3",
   508 => x"124aa3c5",
   509 => x"4aa3c751",
   510 => x"a3c95112",
   511 => x"ce51124a",
   512 => x"51124aa3",
   513 => x"124aa3d0",
   514 => x"4aa3d251",
   515 => x"a3d45112",
   516 => x"d651124a",
   517 => x"51124aa3",
   518 => x"124aa3d8",
   519 => x"4aa3dc51",
   520 => x"a3de5112",
   521 => x"c151124a",
   522 => x"87f8c07e",
   523 => x"99c84974",
   524 => x"87e9c005",
   525 => x"99d04974",
   526 => x"dc87cf05",
   527 => x"87ca0266",
   528 => x"66dc4973",
   529 => x"0298700f",
   530 => x"056e87d3",
   531 => x"c287c6c0",
   532 => x"c048d4c9",
   533 => x"c3e4c050",
   534 => x"e1c248bf",
   535 => x"e1c9c287",
   536 => x"7e50c048",
   537 => x"bfd0c9c2",
   538 => x"c0c1c249",
   539 => x"aa714abf",
   540 => x"87f9fb04",
   541 => x"bff1cdc2",
   542 => x"87c8c005",
   543 => x"bfccc9c2",
   544 => x"87f8c102",
   545 => x"bffcc0c2",
   546 => x"87d8f049",
   547 => x"c1c24970",
   548 => x"a6c459c0",
   549 => x"fcc0c248",
   550 => x"c9c278bf",
   551 => x"c002bfcc",
   552 => x"66c487d8",
   553 => x"ffffcf49",
   554 => x"a999f8ff",
   555 => x"87c5c002",
   556 => x"e1c04cc0",
   557 => x"c04cc187",
   558 => x"66c487dc",
   559 => x"f8ffcf49",
   560 => x"c002a999",
   561 => x"a6c887c8",
   562 => x"c078c048",
   563 => x"a6c887c5",
   564 => x"c878c148",
   565 => x"9c744c66",
   566 => x"87e0c005",
   567 => x"c24966c4",
   568 => x"c4c9c289",
   569 => x"c2914abf",
   570 => x"4abfddcd",
   571 => x"48f8c0c2",
   572 => x"c278a172",
   573 => x"c048c0c1",
   574 => x"87e1f978",
   575 => x"8ef448c0",
   576 => x"0087d9ee",
   577 => x"ff000000",
   578 => x"13ffffff",
   579 => x"1c000009",
   580 => x"46000009",
   581 => x"32335441",
   582 => x"00202020",
   583 => x"31544146",
   584 => x"20202036",
   585 => x"d4ff1e00",
   586 => x"78ffc348",
   587 => x"4f264868",
   588 => x"48d4ff1e",
   589 => x"ff78ffc3",
   590 => x"e1c048d0",
   591 => x"48d4ff78",
   592 => x"cdc278d4",
   593 => x"d4ff48f5",
   594 => x"4f2650bf",
   595 => x"48d0ff1e",
   596 => x"2678e0c0",
   597 => x"ccff1e4f",
   598 => x"99497087",
   599 => x"c087c602",
   600 => x"f105a9fb",
   601 => x"26487187",
   602 => x"5b5e0e4f",
   603 => x"4b710e5c",
   604 => x"f0fe4cc0",
   605 => x"99497087",
   606 => x"87f9c002",
   607 => x"02a9ecc0",
   608 => x"c087f2c0",
   609 => x"c002a9fb",
   610 => x"66cc87eb",
   611 => x"c703acb7",
   612 => x"0266d087",
   613 => x"537187c2",
   614 => x"c2029971",
   615 => x"fe84c187",
   616 => x"497087c3",
   617 => x"87cd0299",
   618 => x"02a9ecc0",
   619 => x"fbc087c7",
   620 => x"d5ff05a9",
   621 => x"0266d087",
   622 => x"97c087c3",
   623 => x"a9ecc07b",
   624 => x"7487c405",
   625 => x"7487c54a",
   626 => x"8a0ac04a",
   627 => x"87c24872",
   628 => x"4c264d26",
   629 => x"4f264b26",
   630 => x"87c9fd1e",
   631 => x"c04a4970",
   632 => x"c904aaf0",
   633 => x"aaf9c087",
   634 => x"c087c301",
   635 => x"c1c18af0",
   636 => x"87c904aa",
   637 => x"01aadac1",
   638 => x"f7c087c3",
   639 => x"2648728a",
   640 => x"5b5e0e4f",
   641 => x"4a710e5c",
   642 => x"724bd4ff",
   643 => x"87e7c049",
   644 => x"029c4c70",
   645 => x"8cc187c2",
   646 => x"c548d0ff",
   647 => x"7bd5c178",
   648 => x"31c64974",
   649 => x"97f7d2c1",
   650 => x"71484abf",
   651 => x"ff7b70b0",
   652 => x"78c448d0",
   653 => x"0e87dbfe",
   654 => x"5d5c5b5e",
   655 => x"7186f80e",
   656 => x"fb7ec04c",
   657 => x"4bc087ea",
   658 => x"97e4ebc0",
   659 => x"a9c049bf",
   660 => x"fb87cf04",
   661 => x"83c187ff",
   662 => x"97e4ebc0",
   663 => x"06ab49bf",
   664 => x"ebc087f1",
   665 => x"02bf97e4",
   666 => x"f8fa87cf",
   667 => x"99497087",
   668 => x"c087c602",
   669 => x"f105a9ec",
   670 => x"fa4bc087",
   671 => x"4d7087e7",
   672 => x"c887e2fa",
   673 => x"dcfa58a6",
   674 => x"c14a7087",
   675 => x"49a4c883",
   676 => x"ad496997",
   677 => x"c087c702",
   678 => x"c005adff",
   679 => x"a4c987e7",
   680 => x"49699749",
   681 => x"02a966c4",
   682 => x"c04887c7",
   683 => x"d405a8ff",
   684 => x"49a4ca87",
   685 => x"aa496997",
   686 => x"c087c602",
   687 => x"c405aaff",
   688 => x"d07ec187",
   689 => x"adecc087",
   690 => x"c087c602",
   691 => x"c405adfb",
   692 => x"c14bc087",
   693 => x"fe026e7e",
   694 => x"eff987e1",
   695 => x"f8487387",
   696 => x"87ecfb8e",
   697 => x"5b5e0e00",
   698 => x"f80e5d5c",
   699 => x"ff4d7186",
   700 => x"1e754bd4",
   701 => x"49facdc2",
   702 => x"c487dbe8",
   703 => x"02987086",
   704 => x"c487ccc4",
   705 => x"d2c148a6",
   706 => x"7578bff9",
   707 => x"87f1fb49",
   708 => x"c548d0ff",
   709 => x"7bd6c178",
   710 => x"a2754ac0",
   711 => x"c17b1149",
   712 => x"aab7cb82",
   713 => x"cc87f304",
   714 => x"7bffc34a",
   715 => x"e0c082c1",
   716 => x"f404aab7",
   717 => x"48d0ff87",
   718 => x"ffc378c4",
   719 => x"c178c57b",
   720 => x"7bc17bd3",
   721 => x"486678c4",
   722 => x"06a8b7c0",
   723 => x"c287f0c2",
   724 => x"4cbfc2ce",
   725 => x"744866c4",
   726 => x"58a6c888",
   727 => x"c1029c74",
   728 => x"c1c287f9",
   729 => x"c0c87ec4",
   730 => x"b7c08c4d",
   731 => x"87c603ac",
   732 => x"4da4c0c8",
   733 => x"cdc24cc0",
   734 => x"49bf97f5",
   735 => x"d10299d0",
   736 => x"c21ec087",
   737 => x"ea49facd",
   738 => x"86c487ff",
   739 => x"c04a4970",
   740 => x"c1c287ee",
   741 => x"cdc21ec4",
   742 => x"ecea49fa",
   743 => x"7086c487",
   744 => x"d0ff4a49",
   745 => x"78c5c848",
   746 => x"6e7bd4c1",
   747 => x"6e7bbf97",
   748 => x"7080c148",
   749 => x"058dc17e",
   750 => x"ff87f0ff",
   751 => x"78c448d0",
   752 => x"c5059a72",
   753 => x"c148c087",
   754 => x"1ec187c7",
   755 => x"49facdc2",
   756 => x"c487dce8",
   757 => x"059c7486",
   758 => x"c487c7fe",
   759 => x"b7c04866",
   760 => x"87d106a8",
   761 => x"48facdc2",
   762 => x"80d078c0",
   763 => x"80f478c0",
   764 => x"bfc6cec2",
   765 => x"4866c478",
   766 => x"01a8b7c0",
   767 => x"ff87d0fd",
   768 => x"78c548d0",
   769 => x"c07bd3c1",
   770 => x"c178c47b",
   771 => x"c087c248",
   772 => x"268ef848",
   773 => x"264c264d",
   774 => x"0e4f264b",
   775 => x"5d5c5b5e",
   776 => x"4b711e0e",
   777 => x"ab4d4cc0",
   778 => x"87e8c004",
   779 => x"1ef7e8c0",
   780 => x"c4029d75",
   781 => x"c24ac087",
   782 => x"724ac187",
   783 => x"87eeeb49",
   784 => x"7e7086c4",
   785 => x"056e84c1",
   786 => x"4c7387c2",
   787 => x"ac7385c1",
   788 => x"87d8ff06",
   789 => x"fe26486e",
   790 => x"711e87f9",
   791 => x"0566c44a",
   792 => x"497287c5",
   793 => x"2687fef9",
   794 => x"5b5e0e4f",
   795 => x"1e0e5d5c",
   796 => x"de494c71",
   797 => x"e2cec291",
   798 => x"9785714d",
   799 => x"ddc1026d",
   800 => x"cecec287",
   801 => x"82744abf",
   802 => x"cefe4972",
   803 => x"487e7087",
   804 => x"f2c00298",
   805 => x"d6cec287",
   806 => x"cb4a704b",
   807 => x"c6d0ff49",
   808 => x"cb4b7487",
   809 => x"cbd3c193",
   810 => x"c083c483",
   811 => x"747be2f3",
   812 => x"dffec049",
   813 => x"c17b7587",
   814 => x"bf97f8d2",
   815 => x"cec21e49",
   816 => x"d5fe49d6",
   817 => x"7486c487",
   818 => x"c7fec049",
   819 => x"c049c087",
   820 => x"c287e6ff",
   821 => x"c048f6cd",
   822 => x"de49c178",
   823 => x"fc2687dc",
   824 => x"6f4c87f1",
   825 => x"6e696461",
   826 => x"2e2e2e67",
   827 => x"5b5e0e00",
   828 => x"4b710e5c",
   829 => x"cecec24a",
   830 => x"497282bf",
   831 => x"7087dcfc",
   832 => x"c4029c4c",
   833 => x"ede74987",
   834 => x"cecec287",
   835 => x"c178c048",
   836 => x"87e6dd49",
   837 => x"0e87fefb",
   838 => x"5d5c5b5e",
   839 => x"c286f40e",
   840 => x"c04dc4c1",
   841 => x"48a6c44c",
   842 => x"cec278c0",
   843 => x"c049bfce",
   844 => x"c1c106a9",
   845 => x"c4c1c287",
   846 => x"c0029848",
   847 => x"e8c087f8",
   848 => x"66c81ef7",
   849 => x"c487c702",
   850 => x"78c048a6",
   851 => x"a6c487c5",
   852 => x"c478c148",
   853 => x"d5e74966",
   854 => x"7086c487",
   855 => x"c484c14d",
   856 => x"80c14866",
   857 => x"c258a6c8",
   858 => x"49bfcece",
   859 => x"87c603ac",
   860 => x"ff059d75",
   861 => x"4cc087c8",
   862 => x"c3029d75",
   863 => x"e8c087e0",
   864 => x"66c81ef7",
   865 => x"cc87c702",
   866 => x"78c048a6",
   867 => x"a6cc87c5",
   868 => x"cc78c148",
   869 => x"d5e64966",
   870 => x"7086c487",
   871 => x"0298487e",
   872 => x"4987e8c2",
   873 => x"699781cb",
   874 => x"0299d049",
   875 => x"c087d6c1",
   876 => x"744aedf3",
   877 => x"c191cb49",
   878 => x"7281cbd3",
   879 => x"c381c879",
   880 => x"497451ff",
   881 => x"cec291de",
   882 => x"85714de2",
   883 => x"7d97c1c2",
   884 => x"c049a5c1",
   885 => x"c9c251e0",
   886 => x"02bf97d4",
   887 => x"84c187d2",
   888 => x"c24ba5c2",
   889 => x"db4ad4c9",
   890 => x"facaff49",
   891 => x"87dbc187",
   892 => x"c049a5cd",
   893 => x"c284c151",
   894 => x"4a6e4ba5",
   895 => x"caff49cb",
   896 => x"c6c187e5",
   897 => x"e9f1c087",
   898 => x"cb49744a",
   899 => x"cbd3c191",
   900 => x"c2797281",
   901 => x"bf97d4c9",
   902 => x"7487d802",
   903 => x"c191de49",
   904 => x"e2cec284",
   905 => x"c283714b",
   906 => x"dd4ad4c9",
   907 => x"f6c9ff49",
   908 => x"7487d887",
   909 => x"c293de4b",
   910 => x"cb83e2ce",
   911 => x"51c049a3",
   912 => x"6e7384c1",
   913 => x"ff49cb4a",
   914 => x"c487dcc9",
   915 => x"80c14866",
   916 => x"c758a6c8",
   917 => x"c5c003ac",
   918 => x"fc056e87",
   919 => x"487487e0",
   920 => x"eef68ef4",
   921 => x"1e731e87",
   922 => x"cb494b71",
   923 => x"cbd3c191",
   924 => x"4aa1c881",
   925 => x"48f7d2c1",
   926 => x"a1c95012",
   927 => x"e4ebc04a",
   928 => x"ca501248",
   929 => x"f8d2c181",
   930 => x"c1501148",
   931 => x"bf97f8d2",
   932 => x"49c01e49",
   933 => x"c287c3f7",
   934 => x"de48f6cd",
   935 => x"d749c178",
   936 => x"f52687d8",
   937 => x"711e87f1",
   938 => x"91cb494a",
   939 => x"81cbd3c1",
   940 => x"481181c8",
   941 => x"58facdc2",
   942 => x"48cecec2",
   943 => x"49c178c0",
   944 => x"2687f7d6",
   945 => x"49c01e4f",
   946 => x"87edf7c0",
   947 => x"711e4f26",
   948 => x"87d20299",
   949 => x"48e0d4c1",
   950 => x"80f750c0",
   951 => x"40e6fac0",
   952 => x"78c4d3c1",
   953 => x"d4c187ce",
   954 => x"d2c148dc",
   955 => x"80fc78fd",
   956 => x"78c5fbc0",
   957 => x"5e0e4f26",
   958 => x"0e5d5c5b",
   959 => x"4d7186f4",
   960 => x"c191cb49",
   961 => x"c881cbd3",
   962 => x"a1ca4aa1",
   963 => x"48a6c47e",
   964 => x"bffed1c2",
   965 => x"bf976e78",
   966 => x"4866c44b",
   967 => x"4b702873",
   968 => x"cc48124c",
   969 => x"9c7058a6",
   970 => x"81c984c1",
   971 => x"b7496997",
   972 => x"87c204ac",
   973 => x"976e4cc0",
   974 => x"66c84abf",
   975 => x"ff317249",
   976 => x"9966c4b9",
   977 => x"30724874",
   978 => x"71484a70",
   979 => x"c2d2c2b0",
   980 => x"ffe1c058",
   981 => x"d449c087",
   982 => x"497587e0",
   983 => x"87f4f3c0",
   984 => x"eef28ef4",
   985 => x"1e731e87",
   986 => x"fe494b71",
   987 => x"497387c8",
   988 => x"f287c3fe",
   989 => x"731e87e1",
   990 => x"c64b711e",
   991 => x"db024aa3",
   992 => x"028ac187",
   993 => x"028a87d6",
   994 => x"8a87dac1",
   995 => x"87fcc002",
   996 => x"e1c0028a",
   997 => x"cb028a87",
   998 => x"87dbc187",
   999 => x"c5fc49c7",
  1000 => x"87dec187",
  1001 => x"bfcecec2",
  1002 => x"87cbc102",
  1003 => x"c288c148",
  1004 => x"c158d2ce",
  1005 => x"cec287c1",
  1006 => x"c002bfd2",
  1007 => x"cec287f9",
  1008 => x"c148bfce",
  1009 => x"d2cec280",
  1010 => x"87ebc058",
  1011 => x"bfcecec2",
  1012 => x"c289c649",
  1013 => x"c059d2ce",
  1014 => x"da03a9b7",
  1015 => x"cecec287",
  1016 => x"d278c048",
  1017 => x"d2cec287",
  1018 => x"87cb02bf",
  1019 => x"bfcecec2",
  1020 => x"c280c648",
  1021 => x"c058d2ce",
  1022 => x"87fed149",
  1023 => x"f1c04973",
  1024 => x"d2f087d2",
  1025 => x"5b5e0e87",
  1026 => x"ff0e5d5c",
  1027 => x"a6dc86d0",
  1028 => x"48a6c859",
  1029 => x"80c478c0",
  1030 => x"7866c4c1",
  1031 => x"78c180c4",
  1032 => x"78c180c4",
  1033 => x"48d2cec2",
  1034 => x"cdc278c1",
  1035 => x"de48bff6",
  1036 => x"87cb05a8",
  1037 => x"7087e0f3",
  1038 => x"59a6cc49",
  1039 => x"e387facf",
  1040 => x"d0e487ee",
  1041 => x"87dde387",
  1042 => x"fbc04c70",
  1043 => x"fbc102ac",
  1044 => x"0566d887",
  1045 => x"c187edc1",
  1046 => x"c44a66c0",
  1047 => x"727e6a82",
  1048 => x"eed1c11e",
  1049 => x"4966c448",
  1050 => x"204aa1c8",
  1051 => x"05aa7141",
  1052 => x"511087f9",
  1053 => x"c0c14a26",
  1054 => x"f9c04866",
  1055 => x"496a78e5",
  1056 => x"517481c7",
  1057 => x"4966c0c1",
  1058 => x"51c181c8",
  1059 => x"4966c0c1",
  1060 => x"51c081c9",
  1061 => x"4966c0c1",
  1062 => x"51c081ca",
  1063 => x"1ed81ec1",
  1064 => x"81c8496a",
  1065 => x"c887c2e3",
  1066 => x"66c4c186",
  1067 => x"01a8c048",
  1068 => x"a6c887c7",
  1069 => x"ce78c148",
  1070 => x"66c4c187",
  1071 => x"d088c148",
  1072 => x"87c358a6",
  1073 => x"d087cee2",
  1074 => x"78c248a6",
  1075 => x"cd029c74",
  1076 => x"66c887e3",
  1077 => x"66c8c148",
  1078 => x"d8cd03a8",
  1079 => x"48a6dc87",
  1080 => x"80e878c0",
  1081 => x"fce078c0",
  1082 => x"c14c7087",
  1083 => x"c205acd0",
  1084 => x"66c487d8",
  1085 => x"87e0e37e",
  1086 => x"a6c84970",
  1087 => x"87e5e059",
  1088 => x"ecc04c70",
  1089 => x"ecc105ac",
  1090 => x"4966c887",
  1091 => x"c0c191cb",
  1092 => x"a1c48166",
  1093 => x"c84d6a4a",
  1094 => x"66c44aa1",
  1095 => x"e6fac052",
  1096 => x"87c1e079",
  1097 => x"029c4c70",
  1098 => x"fbc087d9",
  1099 => x"87d302ac",
  1100 => x"dfff5574",
  1101 => x"4c7087ef",
  1102 => x"87c7029c",
  1103 => x"05acfbc0",
  1104 => x"c087edff",
  1105 => x"c1c255e0",
  1106 => x"7d97c055",
  1107 => x"6e4966d8",
  1108 => x"87db05a9",
  1109 => x"cc4866c8",
  1110 => x"ca04a866",
  1111 => x"4866c887",
  1112 => x"a6cc80c1",
  1113 => x"cc87c858",
  1114 => x"88c14866",
  1115 => x"ff58a6d0",
  1116 => x"7087f2de",
  1117 => x"acd0c14c",
  1118 => x"d487c805",
  1119 => x"80c14866",
  1120 => x"c158a6d8",
  1121 => x"fd02acd0",
  1122 => x"e0c087e8",
  1123 => x"66d848a6",
  1124 => x"4866c478",
  1125 => x"a866e0c0",
  1126 => x"87ebc905",
  1127 => x"48a6e4c0",
  1128 => x"487478c0",
  1129 => x"7088fbc0",
  1130 => x"0298487e",
  1131 => x"4887edc9",
  1132 => x"7e7088cb",
  1133 => x"c1029848",
  1134 => x"c94887cd",
  1135 => x"487e7088",
  1136 => x"c1c40298",
  1137 => x"88c44887",
  1138 => x"98487e70",
  1139 => x"4887ce02",
  1140 => x"7e7088c1",
  1141 => x"c3029848",
  1142 => x"e1c887ec",
  1143 => x"48a6dc87",
  1144 => x"ff78f0c0",
  1145 => x"7087fedc",
  1146 => x"acecc04c",
  1147 => x"87c4c002",
  1148 => x"5ca6e0c0",
  1149 => x"02acecc0",
  1150 => x"dcff87cd",
  1151 => x"4c7087e7",
  1152 => x"05acecc0",
  1153 => x"c087f3ff",
  1154 => x"c002acec",
  1155 => x"dcff87c4",
  1156 => x"1ec087d3",
  1157 => x"66d01eca",
  1158 => x"c191cb49",
  1159 => x"714866c8",
  1160 => x"58a6cc80",
  1161 => x"c44866c8",
  1162 => x"58a6d080",
  1163 => x"49bf66cc",
  1164 => x"87f5dcff",
  1165 => x"1ede1ec1",
  1166 => x"49bf66d4",
  1167 => x"87e9dcff",
  1168 => x"497086d0",
  1169 => x"c08909c0",
  1170 => x"c059a6ec",
  1171 => x"c04866e8",
  1172 => x"eec006a8",
  1173 => x"66e8c087",
  1174 => x"03a8dd48",
  1175 => x"c487e4c0",
  1176 => x"c049bf66",
  1177 => x"c08166e8",
  1178 => x"e8c051e0",
  1179 => x"81c14966",
  1180 => x"81bf66c4",
  1181 => x"c051c1c2",
  1182 => x"c24966e8",
  1183 => x"bf66c481",
  1184 => x"6e51c081",
  1185 => x"e5f9c048",
  1186 => x"c8496e78",
  1187 => x"5166d081",
  1188 => x"81c9496e",
  1189 => x"6e5166d4",
  1190 => x"dc81ca49",
  1191 => x"66d05166",
  1192 => x"d480c148",
  1193 => x"66c858a6",
  1194 => x"a866cc48",
  1195 => x"87cbc004",
  1196 => x"c14866c8",
  1197 => x"58a6cc80",
  1198 => x"cc87e1c5",
  1199 => x"88c14866",
  1200 => x"c558a6d0",
  1201 => x"dcff87d6",
  1202 => x"497087ce",
  1203 => x"59a6ecc0",
  1204 => x"87c4dcff",
  1205 => x"e0c04970",
  1206 => x"66dc59a6",
  1207 => x"a8ecc048",
  1208 => x"87cac005",
  1209 => x"c048a6dc",
  1210 => x"c07866e8",
  1211 => x"d8ff87c4",
  1212 => x"66c887f3",
  1213 => x"c191cb49",
  1214 => x"714866c0",
  1215 => x"4a7e7080",
  1216 => x"496e82c8",
  1217 => x"e8c081ca",
  1218 => x"66dc5166",
  1219 => x"c081c149",
  1220 => x"c18966e8",
  1221 => x"70307148",
  1222 => x"7189c149",
  1223 => x"d1c27a97",
  1224 => x"c049bffe",
  1225 => x"972966e8",
  1226 => x"71484a6a",
  1227 => x"a6f0c098",
  1228 => x"c4496e58",
  1229 => x"c04d6981",
  1230 => x"c44866e0",
  1231 => x"c002a866",
  1232 => x"a6c487c8",
  1233 => x"c078c048",
  1234 => x"a6c487c5",
  1235 => x"c478c148",
  1236 => x"e0c01e66",
  1237 => x"ff49751e",
  1238 => x"c887ced8",
  1239 => x"c04c7086",
  1240 => x"c106acb7",
  1241 => x"857487d4",
  1242 => x"7449e0c0",
  1243 => x"c14b7589",
  1244 => x"714af7d1",
  1245 => x"87eff4fe",
  1246 => x"e4c085c2",
  1247 => x"80c14866",
  1248 => x"58a6e8c0",
  1249 => x"4966ecc0",
  1250 => x"a97081c1",
  1251 => x"87c8c002",
  1252 => x"c048a6c4",
  1253 => x"87c5c078",
  1254 => x"c148a6c4",
  1255 => x"1e66c478",
  1256 => x"c049a4c2",
  1257 => x"887148e0",
  1258 => x"751e4970",
  1259 => x"f8d6ff49",
  1260 => x"c086c887",
  1261 => x"ff01a8b7",
  1262 => x"e4c087c0",
  1263 => x"d1c00266",
  1264 => x"c9496e87",
  1265 => x"66e4c081",
  1266 => x"c0486e51",
  1267 => x"c078f6fb",
  1268 => x"496e87cc",
  1269 => x"51c281c9",
  1270 => x"fdc0486e",
  1271 => x"66c878e5",
  1272 => x"a866cc48",
  1273 => x"87cbc004",
  1274 => x"c14866c8",
  1275 => x"58a6cc80",
  1276 => x"cc87e9c0",
  1277 => x"88c14866",
  1278 => x"c058a6d0",
  1279 => x"d5ff87de",
  1280 => x"4c7087d3",
  1281 => x"c187d5c0",
  1282 => x"c005acc6",
  1283 => x"66d087c8",
  1284 => x"d480c148",
  1285 => x"d4ff58a6",
  1286 => x"4c7087fb",
  1287 => x"c14866d4",
  1288 => x"58a6d880",
  1289 => x"c0029c74",
  1290 => x"66c887cb",
  1291 => x"66c8c148",
  1292 => x"e8f204a8",
  1293 => x"d3d4ff87",
  1294 => x"4866c887",
  1295 => x"c003a8c7",
  1296 => x"cec287e5",
  1297 => x"78c048d2",
  1298 => x"cb4966c8",
  1299 => x"66c0c191",
  1300 => x"4aa1c481",
  1301 => x"52c04a6a",
  1302 => x"4866c879",
  1303 => x"a6cc80c1",
  1304 => x"04a8c758",
  1305 => x"ff87dbff",
  1306 => x"deff8ed0",
  1307 => x"6f4c87e5",
  1308 => x"2a206461",
  1309 => x"3a00202e",
  1310 => x"731e0020",
  1311 => x"9b4b711e",
  1312 => x"c287c602",
  1313 => x"c048cece",
  1314 => x"c21ec778",
  1315 => x"49bfcece",
  1316 => x"cbd3c11e",
  1317 => x"f6cdc21e",
  1318 => x"e8ed49bf",
  1319 => x"c286cc87",
  1320 => x"49bff6cd",
  1321 => x"7387e7e8",
  1322 => x"87c7029b",
  1323 => x"49cbd3c1",
  1324 => x"ff87f3df",
  1325 => x"0087e0dd",
  1326 => x"00000100",
  1327 => x"45208000",
  1328 => x"00746978",
  1329 => x"61422080",
  1330 => x"69006b63",
  1331 => x"a200000c",
  1332 => x"00000023",
  1333 => x"0c690000",
  1334 => x"23c00000",
  1335 => x"00000000",
  1336 => x"000c6900",
  1337 => x"0023de00",
  1338 => x"00000000",
  1339 => x"00000c69",
  1340 => x"000023fc",
  1341 => x"69000000",
  1342 => x"1a00000c",
  1343 => x"00000024",
  1344 => x"0c690000",
  1345 => x"24380000",
  1346 => x"00000000",
  1347 => x"000c6900",
  1348 => x"00245600",
  1349 => x"00000000",
  1350 => x"00000ea6",
  1351 => x"00000000",
  1352 => x"76000000",
  1353 => x"0000000f",
  1354 => x"00000000",
  1355 => x"fe1e0000",
  1356 => x"78c048f0",
  1357 => x"097909cd",
  1358 => x"1e1e4f26",
  1359 => x"7ebff0fe",
  1360 => x"4f262648",
  1361 => x"48f0fe1e",
  1362 => x"4f2678c1",
  1363 => x"48f0fe1e",
  1364 => x"4f2678c0",
  1365 => x"c04a711e",
  1366 => x"4f265252",
  1367 => x"5c5b5e0e",
  1368 => x"86f40e5d",
  1369 => x"6d974d71",
  1370 => x"4ca5c17e",
  1371 => x"c8486c97",
  1372 => x"486e58a6",
  1373 => x"05a866c4",
  1374 => x"48ff87c5",
  1375 => x"ff87e6c0",
  1376 => x"a5c287ca",
  1377 => x"4b6c9749",
  1378 => x"974ba371",
  1379 => x"6c974b6b",
  1380 => x"c1486e7e",
  1381 => x"58a6c880",
  1382 => x"a6cc98c7",
  1383 => x"7c977058",
  1384 => x"7387e1fe",
  1385 => x"268ef448",
  1386 => x"264c264d",
  1387 => x"0e4f264b",
  1388 => x"0e5c5b5e",
  1389 => x"4c7186f4",
  1390 => x"c34a66d8",
  1391 => x"a4c29aff",
  1392 => x"496c974b",
  1393 => x"7249a173",
  1394 => x"7e6c9751",
  1395 => x"80c1486e",
  1396 => x"c758a6c8",
  1397 => x"58a6cc98",
  1398 => x"8ef45470",
  1399 => x"1e87caff",
  1400 => x"87e8fd1e",
  1401 => x"494abfe0",
  1402 => x"99c0e0c0",
  1403 => x"7287cb02",
  1404 => x"f4d1c21e",
  1405 => x"87f7fe49",
  1406 => x"fdfc86c4",
  1407 => x"fd7e7087",
  1408 => x"262687c2",
  1409 => x"d1c21e4f",
  1410 => x"c7fd49f4",
  1411 => x"dfd7c187",
  1412 => x"87dafc49",
  1413 => x"2687fec2",
  1414 => x"1e731e4f",
  1415 => x"49f4d1c2",
  1416 => x"7087f9fc",
  1417 => x"aab7c04a",
  1418 => x"87ccc204",
  1419 => x"05aaf0c3",
  1420 => x"dbc187c9",
  1421 => x"78c148c4",
  1422 => x"c387edc1",
  1423 => x"c905aae0",
  1424 => x"c8dbc187",
  1425 => x"c178c148",
  1426 => x"dbc187de",
  1427 => x"c602bfc8",
  1428 => x"a2c0c287",
  1429 => x"7287c24b",
  1430 => x"c4dbc14b",
  1431 => x"e0c002bf",
  1432 => x"c4497387",
  1433 => x"c19129b7",
  1434 => x"7381e4dc",
  1435 => x"c29acf4a",
  1436 => x"7248c192",
  1437 => x"ff4a7030",
  1438 => x"694872ba",
  1439 => x"db797098",
  1440 => x"c4497387",
  1441 => x"c19129b7",
  1442 => x"7381e4dc",
  1443 => x"c29acf4a",
  1444 => x"7248c392",
  1445 => x"484a7030",
  1446 => x"7970b069",
  1447 => x"48c8dbc1",
  1448 => x"dbc178c0",
  1449 => x"78c048c4",
  1450 => x"49f4d1c2",
  1451 => x"7087edfa",
  1452 => x"aab7c04a",
  1453 => x"87f4fd03",
  1454 => x"87c448c0",
  1455 => x"4c264d26",
  1456 => x"4f264b26",
  1457 => x"00000000",
  1458 => x"00000000",
  1459 => x"494a711e",
  1460 => x"2687c6fd",
  1461 => x"4ac01e4f",
  1462 => x"91c44972",
  1463 => x"81e4dcc1",
  1464 => x"82c179c0",
  1465 => x"04aab7d0",
  1466 => x"4f2687ee",
  1467 => x"5c5b5e0e",
  1468 => x"4d710e5d",
  1469 => x"7587d5f9",
  1470 => x"2ab7c44a",
  1471 => x"e4dcc192",
  1472 => x"cf4c7582",
  1473 => x"6a94c29c",
  1474 => x"2b744b49",
  1475 => x"48c29bc3",
  1476 => x"4c703074",
  1477 => x"4874bcff",
  1478 => x"7a709871",
  1479 => x"7387e5f8",
  1480 => x"87d8fe48",
  1481 => x"00000000",
  1482 => x"00000000",
  1483 => x"00000000",
  1484 => x"00000000",
  1485 => x"00000000",
  1486 => x"00000000",
  1487 => x"00000000",
  1488 => x"00000000",
  1489 => x"00000000",
  1490 => x"00000000",
  1491 => x"00000000",
  1492 => x"00000000",
  1493 => x"00000000",
  1494 => x"00000000",
  1495 => x"00000000",
  1496 => x"00000000",
  1497 => x"48d0ff1e",
  1498 => x"7178e1c8",
  1499 => x"08d4ff48",
  1500 => x"4866c478",
  1501 => x"7808d4ff",
  1502 => x"711e4f26",
  1503 => x"4966c44a",
  1504 => x"ff49721e",
  1505 => x"d0ff87de",
  1506 => x"78e0c048",
  1507 => x"1e4f2626",
  1508 => x"4b711e73",
  1509 => x"1e4966c8",
  1510 => x"e0c14a73",
  1511 => x"d9ff49a2",
  1512 => x"87c42687",
  1513 => x"4c264d26",
  1514 => x"4f264b26",
  1515 => x"711e731e",
  1516 => x"b7c24b4a",
  1517 => x"87c803ab",
  1518 => x"c34a49a3",
  1519 => x"87c79aff",
  1520 => x"4a49a3ce",
  1521 => x"c89affc3",
  1522 => x"721e4966",
  1523 => x"87eafe49",
  1524 => x"87d4ff26",
  1525 => x"4ad4ff1e",
  1526 => x"ff7affc3",
  1527 => x"e1c048d0",
  1528 => x"c27ade78",
  1529 => x"7abffed1",
  1530 => x"28c84849",
  1531 => x"48717a70",
  1532 => x"7a7028d0",
  1533 => x"28d84871",
  1534 => x"d0ff7a70",
  1535 => x"78e0c048",
  1536 => x"ff1e4f26",
  1537 => x"c9c848d0",
  1538 => x"ff487178",
  1539 => x"267808d4",
  1540 => x"4a711e4f",
  1541 => x"ff87eb49",
  1542 => x"78c848d0",
  1543 => x"731e4f26",
  1544 => x"c24b711e",
  1545 => x"02bfced2",
  1546 => x"ebc287c3",
  1547 => x"48d0ff87",
  1548 => x"7378c9c8",
  1549 => x"b1e0c049",
  1550 => x"7148d4ff",
  1551 => x"c2d2c278",
  1552 => x"c878c048",
  1553 => x"87c50266",
  1554 => x"c249ffc3",
  1555 => x"c249c087",
  1556 => x"cc59cad2",
  1557 => x"87c60266",
  1558 => x"4ad5d5c5",
  1559 => x"ffcf87c4",
  1560 => x"d2c24aff",
  1561 => x"d2c25ace",
  1562 => x"78c148ce",
  1563 => x"4d2687c4",
  1564 => x"4b264c26",
  1565 => x"5e0e4f26",
  1566 => x"0e5d5c5b",
  1567 => x"d2c24a71",
  1568 => x"724cbfca",
  1569 => x"87cb029a",
  1570 => x"c191c849",
  1571 => x"714bd4e0",
  1572 => x"c187c483",
  1573 => x"c04bd4e4",
  1574 => x"7449134d",
  1575 => x"c6d2c299",
  1576 => x"d4ffb9bf",
  1577 => x"c1787148",
  1578 => x"c8852cb7",
  1579 => x"e804adb7",
  1580 => x"c2d2c287",
  1581 => x"80c848bf",
  1582 => x"58c6d2c2",
  1583 => x"1e87effe",
  1584 => x"4b711e73",
  1585 => x"029a4a13",
  1586 => x"497287cb",
  1587 => x"1387e7fe",
  1588 => x"f5059a4a",
  1589 => x"87dafe87",
  1590 => x"c2d2c21e",
  1591 => x"d2c249bf",
  1592 => x"a1c148c2",
  1593 => x"b7c0c478",
  1594 => x"87db03a9",
  1595 => x"c248d4ff",
  1596 => x"78bfc6d2",
  1597 => x"bfc2d2c2",
  1598 => x"c2d2c249",
  1599 => x"78a1c148",
  1600 => x"a9b7c0c4",
  1601 => x"ff87e504",
  1602 => x"78c848d0",
  1603 => x"48ced2c2",
  1604 => x"4f2678c0",
  1605 => x"00000000",
  1606 => x"00000000",
  1607 => x"5f000000",
  1608 => x"0000005f",
  1609 => x"00030300",
  1610 => x"00000303",
  1611 => x"147f7f14",
  1612 => x"00147f7f",
  1613 => x"6b2e2400",
  1614 => x"00123a6b",
  1615 => x"18366a4c",
  1616 => x"0032566c",
  1617 => x"594f7e30",
  1618 => x"40683a77",
  1619 => x"07040000",
  1620 => x"00000003",
  1621 => x"3e1c0000",
  1622 => x"00004163",
  1623 => x"63410000",
  1624 => x"00001c3e",
  1625 => x"1c3e2a08",
  1626 => x"082a3e1c",
  1627 => x"3e080800",
  1628 => x"0008083e",
  1629 => x"e0800000",
  1630 => x"00000060",
  1631 => x"08080800",
  1632 => x"00080808",
  1633 => x"60000000",
  1634 => x"00000060",
  1635 => x"18306040",
  1636 => x"0103060c",
  1637 => x"597f3e00",
  1638 => x"003e7f4d",
  1639 => x"7f060400",
  1640 => x"0000007f",
  1641 => x"71634200",
  1642 => x"00464f59",
  1643 => x"49632200",
  1644 => x"00367f49",
  1645 => x"13161c18",
  1646 => x"00107f7f",
  1647 => x"45672700",
  1648 => x"00397d45",
  1649 => x"4b7e3c00",
  1650 => x"00307949",
  1651 => x"71010100",
  1652 => x"00070f79",
  1653 => x"497f3600",
  1654 => x"00367f49",
  1655 => x"494f0600",
  1656 => x"001e3f69",
  1657 => x"66000000",
  1658 => x"00000066",
  1659 => x"e6800000",
  1660 => x"00000066",
  1661 => x"14080800",
  1662 => x"00222214",
  1663 => x"14141400",
  1664 => x"00141414",
  1665 => x"14222200",
  1666 => x"00080814",
  1667 => x"51030200",
  1668 => x"00060f59",
  1669 => x"5d417f3e",
  1670 => x"001e1f55",
  1671 => x"097f7e00",
  1672 => x"007e7f09",
  1673 => x"497f7f00",
  1674 => x"00367f49",
  1675 => x"633e1c00",
  1676 => x"00414141",
  1677 => x"417f7f00",
  1678 => x"001c3e63",
  1679 => x"497f7f00",
  1680 => x"00414149",
  1681 => x"097f7f00",
  1682 => x"00010109",
  1683 => x"417f3e00",
  1684 => x"007a7b49",
  1685 => x"087f7f00",
  1686 => x"007f7f08",
  1687 => x"7f410000",
  1688 => x"0000417f",
  1689 => x"40602000",
  1690 => x"003f7f40",
  1691 => x"1c087f7f",
  1692 => x"00416336",
  1693 => x"407f7f00",
  1694 => x"00404040",
  1695 => x"0c067f7f",
  1696 => x"007f7f06",
  1697 => x"0c067f7f",
  1698 => x"007f7f18",
  1699 => x"417f3e00",
  1700 => x"003e7f41",
  1701 => x"097f7f00",
  1702 => x"00060f09",
  1703 => x"61417f3e",
  1704 => x"00407e7f",
  1705 => x"097f7f00",
  1706 => x"00667f19",
  1707 => x"4d6f2600",
  1708 => x"00327b59",
  1709 => x"7f010100",
  1710 => x"0001017f",
  1711 => x"407f3f00",
  1712 => x"003f7f40",
  1713 => x"703f0f00",
  1714 => x"000f3f70",
  1715 => x"18307f7f",
  1716 => x"007f7f30",
  1717 => x"1c366341",
  1718 => x"4163361c",
  1719 => x"7c060301",
  1720 => x"0103067c",
  1721 => x"4d597161",
  1722 => x"00414347",
  1723 => x"7f7f0000",
  1724 => x"00004141",
  1725 => x"0c060301",
  1726 => x"40603018",
  1727 => x"41410000",
  1728 => x"00007f7f",
  1729 => x"03060c08",
  1730 => x"00080c06",
  1731 => x"80808080",
  1732 => x"00808080",
  1733 => x"03000000",
  1734 => x"00000407",
  1735 => x"54742000",
  1736 => x"00787c54",
  1737 => x"447f7f00",
  1738 => x"00387c44",
  1739 => x"447c3800",
  1740 => x"00004444",
  1741 => x"447c3800",
  1742 => x"007f7f44",
  1743 => x"547c3800",
  1744 => x"00185c54",
  1745 => x"7f7e0400",
  1746 => x"00000505",
  1747 => x"a4bc1800",
  1748 => x"007cfca4",
  1749 => x"047f7f00",
  1750 => x"00787c04",
  1751 => x"3d000000",
  1752 => x"0000407d",
  1753 => x"80808000",
  1754 => x"00007dfd",
  1755 => x"107f7f00",
  1756 => x"00446c38",
  1757 => x"3f000000",
  1758 => x"0000407f",
  1759 => x"180c7c7c",
  1760 => x"00787c0c",
  1761 => x"047c7c00",
  1762 => x"00787c04",
  1763 => x"447c3800",
  1764 => x"00387c44",
  1765 => x"24fcfc00",
  1766 => x"00183c24",
  1767 => x"243c1800",
  1768 => x"00fcfc24",
  1769 => x"047c7c00",
  1770 => x"00080c04",
  1771 => x"545c4800",
  1772 => x"00207454",
  1773 => x"7f3f0400",
  1774 => x"00004444",
  1775 => x"407c3c00",
  1776 => x"007c7c40",
  1777 => x"603c1c00",
  1778 => x"001c3c60",
  1779 => x"30607c3c",
  1780 => x"003c7c60",
  1781 => x"10386c44",
  1782 => x"00446c38",
  1783 => x"e0bc1c00",
  1784 => x"001c3c60",
  1785 => x"74644400",
  1786 => x"00444c5c",
  1787 => x"3e080800",
  1788 => x"00414177",
  1789 => x"7f000000",
  1790 => x"0000007f",
  1791 => x"77414100",
  1792 => x"0008083e",
  1793 => x"03010102",
  1794 => x"00010202",
  1795 => x"7f7f7f7f",
  1796 => x"007f7f7f",
  1797 => x"1c1c0808",
  1798 => x"7f7f3e3e",
  1799 => x"3e3e7f7f",
  1800 => x"08081c1c",
  1801 => x"7c181000",
  1802 => x"0010187c",
  1803 => x"7c301000",
  1804 => x"0010307c",
  1805 => x"60603010",
  1806 => x"00061e78",
  1807 => x"183c6642",
  1808 => x"0042663c",
  1809 => x"c26a3878",
  1810 => x"00386cc6",
  1811 => x"60000060",
  1812 => x"00600000",
  1813 => x"5c5b5e0e",
  1814 => x"711e0e5d",
  1815 => x"dfd2c24c",
  1816 => x"4bc04dbf",
  1817 => x"ab741ec0",
  1818 => x"c487c702",
  1819 => x"78c048a6",
  1820 => x"a6c487c5",
  1821 => x"c478c148",
  1822 => x"49731e66",
  1823 => x"c887dfee",
  1824 => x"49e0c086",
  1825 => x"c487efef",
  1826 => x"496a4aa5",
  1827 => x"f187f0f0",
  1828 => x"85cb87c6",
  1829 => x"b7c883c1",
  1830 => x"c7ff04ab",
  1831 => x"4d262687",
  1832 => x"4b264c26",
  1833 => x"711e4f26",
  1834 => x"e3d2c24a",
  1835 => x"e3d2c25a",
  1836 => x"4978c748",
  1837 => x"2687ddfe",
  1838 => x"1e731e4f",
  1839 => x"b7c04a71",
  1840 => x"87d303aa",
  1841 => x"bfe6ffc1",
  1842 => x"c187c405",
  1843 => x"c087c24b",
  1844 => x"eaffc14b",
  1845 => x"c187c45b",
  1846 => x"c15aeaff",
  1847 => x"4abfe6ff",
  1848 => x"c0c19ac1",
  1849 => x"e8ec49a2",
  1850 => x"c148fc87",
  1851 => x"78bfe6ff",
  1852 => x"1e87effe",
  1853 => x"66c44a71",
  1854 => x"ea49721e",
  1855 => x"262687ee",
  1856 => x"4a711e4f",
  1857 => x"c348d4ff",
  1858 => x"d0ff78ff",
  1859 => x"78e1c048",
  1860 => x"c148d4ff",
  1861 => x"c4497278",
  1862 => x"ff787131",
  1863 => x"e0c048d0",
  1864 => x"1e4f2678",
  1865 => x"bfe6ffc1",
  1866 => x"87e0e649",
  1867 => x"48d7d2c2",
  1868 => x"c278bfe8",
  1869 => x"ec48d3d2",
  1870 => x"d2c278bf",
  1871 => x"494abfd7",
  1872 => x"c899ffc3",
  1873 => x"48722ab7",
  1874 => x"d2c2b071",
  1875 => x"4f2658df",
  1876 => x"5c5b5e0e",
  1877 => x"4b710e5d",
  1878 => x"c287c8ff",
  1879 => x"c048d2d2",
  1880 => x"e6497350",
  1881 => x"497087c6",
  1882 => x"cb9cc24c",
  1883 => x"fdc949ee",
  1884 => x"4d497087",
  1885 => x"97d2d2c2",
  1886 => x"e2c105bf",
  1887 => x"4966d087",
  1888 => x"bfdbd2c2",
  1889 => x"87d60599",
  1890 => x"c24966d4",
  1891 => x"99bfd3d2",
  1892 => x"7387cb05",
  1893 => x"87d4e549",
  1894 => x"c1029870",
  1895 => x"4cc187c1",
  1896 => x"7587c0fe",
  1897 => x"87d2c949",
  1898 => x"c6029870",
  1899 => x"d2d2c287",
  1900 => x"c250c148",
  1901 => x"bf97d2d2",
  1902 => x"87e3c005",
  1903 => x"bfdbd2c2",
  1904 => x"9966d049",
  1905 => x"87d6ff05",
  1906 => x"bfd3d2c2",
  1907 => x"9966d449",
  1908 => x"87caff05",
  1909 => x"d3e44973",
  1910 => x"05987087",
  1911 => x"7487fffe",
  1912 => x"87fafa48",
  1913 => x"5c5b5e0e",
  1914 => x"86f80e5d",
  1915 => x"ec4c4dc0",
  1916 => x"a6c47ebf",
  1917 => x"dfd2c248",
  1918 => x"1ec178bf",
  1919 => x"49c71ec0",
  1920 => x"c887cdfd",
  1921 => x"02987086",
  1922 => x"49ff87cd",
  1923 => x"c187eafa",
  1924 => x"d7e349da",
  1925 => x"c24dc187",
  1926 => x"bf97d2d2",
  1927 => x"c187cf02",
  1928 => x"49bfdeff",
  1929 => x"ffc1b9c1",
  1930 => x"fb7159e2",
  1931 => x"d2c287d3",
  1932 => x"c14bbfd7",
  1933 => x"05bfe6ff",
  1934 => x"c387e9c0",
  1935 => x"ebe249fd",
  1936 => x"49fac387",
  1937 => x"7387e5e2",
  1938 => x"99ffc349",
  1939 => x"49c01e71",
  1940 => x"7387e0fa",
  1941 => x"29b7c849",
  1942 => x"49c11e71",
  1943 => x"c887d4fa",
  1944 => x"87f5c586",
  1945 => x"bfdbd2c2",
  1946 => x"dd029b4b",
  1947 => x"e2ffc187",
  1948 => x"c5c649bf",
  1949 => x"05987087",
  1950 => x"4bc087c4",
  1951 => x"e0c287d2",
  1952 => x"87eac549",
  1953 => x"58e6ffc1",
  1954 => x"ffc187c6",
  1955 => x"78c048e2",
  1956 => x"99c24973",
  1957 => x"c387cd05",
  1958 => x"cfe149eb",
  1959 => x"c2497087",
  1960 => x"87c20299",
  1961 => x"49734cfb",
  1962 => x"cd0599c1",
  1963 => x"49f4c387",
  1964 => x"7087f9e0",
  1965 => x"0299c249",
  1966 => x"4cfa87c2",
  1967 => x"99c84973",
  1968 => x"c387cd05",
  1969 => x"e3e049f5",
  1970 => x"c2497087",
  1971 => x"87d50299",
  1972 => x"bfe3d2c2",
  1973 => x"4887ca02",
  1974 => x"d2c288c1",
  1975 => x"c2c058e7",
  1976 => x"c14cff87",
  1977 => x"c449734d",
  1978 => x"87ce0599",
  1979 => x"ff49f2c3",
  1980 => x"7087f9df",
  1981 => x"0299c249",
  1982 => x"d2c287dc",
  1983 => x"487ebfe3",
  1984 => x"03a8b7c7",
  1985 => x"6e87cbc0",
  1986 => x"c280c148",
  1987 => x"c058e7d2",
  1988 => x"4cfe87c2",
  1989 => x"fdc34dc1",
  1990 => x"cfdfff49",
  1991 => x"c2497087",
  1992 => x"87d50299",
  1993 => x"bfe3d2c2",
  1994 => x"87c9c002",
  1995 => x"48e3d2c2",
  1996 => x"c2c078c0",
  1997 => x"c14cfd87",
  1998 => x"49fac34d",
  1999 => x"87ecdeff",
  2000 => x"99c24970",
  2001 => x"87d9c002",
  2002 => x"bfe3d2c2",
  2003 => x"a8b7c748",
  2004 => x"87c9c003",
  2005 => x"48e3d2c2",
  2006 => x"c2c078c7",
  2007 => x"c14cfc87",
  2008 => x"acb7c04d",
  2009 => x"87d3c003",
  2010 => x"c14866c4",
  2011 => x"7e7080d8",
  2012 => x"c002bf6e",
  2013 => x"744b87c5",
  2014 => x"c00f7349",
  2015 => x"1ef0c31e",
  2016 => x"f749dac1",
  2017 => x"86c887ca",
  2018 => x"c0029870",
  2019 => x"d2c287d8",
  2020 => x"6e7ebfe3",
  2021 => x"c491cb49",
  2022 => x"82714a66",
  2023 => x"c5c0026a",
  2024 => x"496e4b87",
  2025 => x"9d750f73",
  2026 => x"87c8c002",
  2027 => x"bfe3d2c2",
  2028 => x"87e0f249",
  2029 => x"bfeaffc1",
  2030 => x"87ddc002",
  2031 => x"87fac049",
  2032 => x"c0029870",
  2033 => x"d2c287d3",
  2034 => x"f249bfe3",
  2035 => x"49c087c6",
  2036 => x"c187e6f3",
  2037 => x"c048eaff",
  2038 => x"f38ef878",
  2039 => x"000087c0",
  2040 => x"00000000",
  2041 => x"00000000",
  2042 => x"00000000",
  2043 => x"711e0000",
  2044 => x"bfc8ff4a",
  2045 => x"48a17249",
  2046 => x"ff1e4f26",
  2047 => x"fe89bfc8",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
